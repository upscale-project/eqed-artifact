
module dff(
input wire d,
output wire q);

assign q = ~d;
endmodule
