module spc_eqed (


spc spc0(
  .vnw_ary0                 (SPC_VNW[ 0 ]),
  .vnw_ary1		    (SPC_VNW[ 0 ]),
  .gclk				  ( cmp_gclk_c3_spc0 ), // cmp_gclk_c1_r[1]) ,
  .tcu_clk_stop ( gl_spc0_clk_stop ),	// staged clk_stop
  .cpx_spc_data_cx	    (cpx_spc0_data_cx2[ 145 : 0 ]	 ),// sparc core
  .pcx_spc_grant_px	    (pcx_spc0_grant_px[ 8 : 0 ]	 ),
  .spc_pcx_req_pq	    (spc0_pcx_req_pq[ 8 : 0 ]	 ),
  .spc_pcx_atm_pq	    (spc0_pcx_atm_pq[ 8 : 0 ]	 ),
  .spc_pcx_data_pa	    (spc0_pcx_data_pa[ 129 : 0 ]	 ),
  .spc_hardstop_request	    (spc0_hardstop_request),
  .spc_softstop_request	    (spc0_softstop_request),
  .spc_trigger_pulse	    (spc0_trigger_pulse),
  .tcu_ss_mode		    (tcu_ss_mode[ 0 ]),
  .tcu_do_mode		    (tcu_do_mode[ 0 ]),
  .tcu_ss_request	    (tcu_ss_request_t1lff_0),
  .spc_ss_complete	    (spc0_ss_complete),
  .tcu_aclk		    (tcu_spc0_aclk		 ),
  .tcu_bclk		    (tcu_spc0_bclk		 ),
  .tcu_scan_en		    (tcu_spc0_scan_en		 ),
  .tcu_se_scancollar_in	    (tcu_spc0_se_scancollar_in	 ),
  .tcu_se_scancollar_out    (tcu_spc0_se_scancollar_out	 ),
  .tcu_array_wr_inhibit	    (tcu_spc0_array_wr_inhibit	 ),
  .tcu_core_running	    (ncu_spc0_core_running[ 7 : 0 ]	 ),
  .spc_core_running_status  (spc0_ncu_core_running_status[ 7 : 0 ]),
  .const_cpuid		    ({1'b0, 1'b0, 1'b0}		 ),//No 3'b101 to Astro.
  .power_throttle	    (mio_spc_pwr_throttle_0[ 2 : 0 ]),
  .scan_out		    (spc0_tcu_scan_in[ 1 : 0 ]	 ),
  .scan_in		    (tcu_spc0_scan_out[ 1 : 0 ]	 ),
  .spc_dbg_instr_cmt_grp0   (spc0_dbg0_instr_cmt_grp0[ 1 : 0 ]),
  .spc_dbg_instr_cmt_grp1   (spc0_dbg0_instr_cmt_grp1[ 1 : 0 ]),
  .tcu_spc_mbist_start	    (tcu_spc0_mbist_start_t1lff_0),
  .spc_mbist_done	    (spc0_tcu_mbist_done    ),
  .spc_mbist_fail	    (spc0_tcu_mbist_fail    ),
  .tcu_spc_mbist_scan_in    (tcu_spc0_mbist_scan_in	 ),
  .spc_tcu_mbist_scan_out   (spc0_tcu_mbist_scan_out	 ),
  .dmo_din		    (36'b0			 ),
  .dmo_dout		    (spc0_dmo_dout[ 35 : 0 ]	 ),
  .dmo_coresel		    (1'b0			 ),
  .tcu_spc_lbist_start	    (tcu_spc_lbist_start[ 0 ]	 ),
  .tcu_spc_lbist_scan_in    (tcu_spc_lbist_scan_in[ 0 ]	 ),
  .spc_tcu_lbist_done	    (spc0_tcu_lbist_done	 ),
  .spc_tcu_lbist_scan_out   (spc0_tcu_lbist_scan_out	 ),
  .tcu_shscan_pce_ov	    (tcu_spc_shscan_pce_ov	 ),
  .tcu_shscan_aclk	    (tcu_spc_shscan_aclk	 ),
  .tcu_shscan_bclk	    (tcu_spc_shscan_bclk	 ),
  .tcu_shscan_scan_en	    (tcu_spc_shscan_scan_en	 ),
  .tcu_shscanid		    (tcu_spc_shscanid[ 2 : 0 ]	 ),
  .tcu_shscan_scan_in	    (tcu_spc0_shscan_scan_out	 ),
  .spc_shscan_scan_out	    (spc0_tcu_shscan_scan_in	 ),
  .tcu_shscan_clk_stop	    (tcu_spc0_shscan_clk_stop	 ),
  .efu_spc_fuse_data	    (efu_spc0246_fuse_data	 ),
  .efu_spc_fuse_ixfer_en    (efu_spc0_fuse_ixfer_en	 ),
  .efu_spc_fuse_iclr	    (efu_spc0_fuse_iclr		 ),
  .efu_spc_fuse_dxfer_en    (efu_spc0_fuse_dxfer_en	 ),
  .efu_spc_fuse_dclr	    (efu_spc0_fuse_dclr		 ),
  .spc_efu_fuse_dxfer_en    (spc0_efu_fuse_dxfer_en	 ),
  .spc_efu_fuse_ixfer_en    (spc0_efu_fuse_ixfer_en	 ),
  .spc_efu_fuse_ddata	    (spc0_efu_fuse_ddata	 ),
  .spc_efu_fuse_idata	    (spc0_efu_fuse_idata	 ),
  .ccu_slow_cmp_sync_en ( gl_io_cmp_sync_en_c3t0 ),	// gl_io_cmp_sync_en_c3t  - for int6.1
  .ccu_cmp_slow_sync_en ( gl_cmp_io_sync_en_c3t0 ),	// gl_cmp_io_sync_en_c3t  - for int6.1
  .hver_mask_minor_rev	    (spc_revid_out[ 3 : 0 ]        ),
  .tcu_pce_ov(tcu_pce_ov),
  .tcu_dectest(tcu_dectest),
  .tcu_muxtest(tcu_muxtest),
  .rst_wmr_protect(rst_wmr_protect),
  .cluster_arst_l(cluster_arst_l),
  .tcu_mbist_bisi_en(tcu_mbist_bisi_en),
  .tcu_mbist_user_mode(tcu_mbist_user_mode),
  .ncu_cmp_tick_enable(ncu_cmp_tick_enable),
  .ncu_wmr_vec_mask(ncu_wmr_vec_mask),
  .ncu_spc_pm(ncu_spc_pm),
  .ncu_spc_ba01(ncu_spc_ba01),
  .ncu_spc_ba23(ncu_spc_ba23),
  .ncu_spc_ba45(ncu_spc_ba45),
  .ncu_spc_ba67(ncu_spc_ba67),
  .tcu_spc_lbist_pgm(tcu_spc_lbist_pgm),
  .tcu_spc_test_mode(tcu_spc0_test_mode),
  .dmo_icmuxctl(dmo_icmuxctl),
  .dmo_dcmuxctl(dmo_dcmuxctl),
  .tcu_atpg_mode(tcu_atpg_mode),
  .ncu_spc_l2_idx_hash_en(ncu_spc_l2_idx_hash_en)
            );

i














































l2t l2t0(
.l2t_lstg_in		    ({
                              148'b0,
			      l2t1_mcu0_rd_req,
			      l2t1_mcu0_rd_dummy_req,
			      l2t1_mcu0_rd_req_id[ 2 : 0 ],
			      l2t1_mcu0_wr_req,
			      l2t1_mcu0_addr_5,
			      l2t1_mcu0_addr[ 39 : 31 ],
			      4'b0,
			      l2t1_mcu0_addr[ 30 : 7 ]}
                            ),
  .l2t_lstg_out		    ({
                              unconnectedt0lff[ 191 : 44 ],
			      l2t1_mcu0_rd_req_t0lff,
			      l2t1_mcu0_rd_dummy_req_t0lff,
			      l2t1_mcu0_rd_req_id_t0lff[ 2 : 0 ],
			      l2t1_mcu0_wr_req_t0lff,
			      l2t1_mcu0_addr_5_t0lff,
			      l2t1_mcu0_addr_t0lff[ 39 : 31 ],
			      unconnectedt0lff[ 27 : 24 ],
			      l2t1_mcu0_addr_t0lff[ 30 : 7 ]}
                            ),
//  .l2t_lstg_in		    (192'b0),
//  .l2t_lstg_out		    (unconnectedt0lff[191:0]),
//  .l2t_rstg_in		    (192'b0),
//  .l2t_rstg_out		    (unconnectedt0rff[191:0]),
  .l2t_rstg_in       	    ({111'b0,
                             l2b0_sio_parity[ 1 : 0 ],
                             79'b0
                             }
                            ),
  .l2t_rstg_out		    ({unconnectedt0rff[ 191 : 81 ],
                             l2b0_sio_parity_t0rff[ 1 : 0 ],
                             unconnectedt0rff[ 78 : 0 ]
                             }
                            ),
  .l2t_siu_delay	    (1'b0),
  .l2t_tcu_dmo_out_prev     (39'b0                       ), 
  .l2t_tcu_dmo_out          (l2t0_dmo_dout[ 38 : 0 ]         ),
  .tcu_l2t_coresel          (1'b0                        ),
  .tcu_l2t_tag_or_data_sel  (dmo_tagmuxctl               ),
  .ccu_slow_cmp_sync_en ( gl_io_cmp_sync_en_c3t ),
  .ccu_cmp_slow_sync_en ( gl_cmp_io_sync_en_c3t ),
  .l2t_dbg_sii_iq_dequeue   (l2t0_dbg0_sii_iq_dequeue	 ),
  .l2t_dbg_sii_wib_dequeue  (l2t0_dbg0_sii_wib_dequeue 	 ),
  .l2t_dbg_xbar_vcid	    (l2t0_dbg0_xbar_vcid[ 5 : 0 ]	 ),
  .l2t_dbg_err_event	    (l2t0_dbg0_err_event		 ),
  .l2t_dbg_pa_match	    (l2t0_dbg0_pa_match		 ),
  .l2t_cpx_req_cq           (sctag0_cpx_req_cq[ 7 : 0 ]      ),// sctag
  .l2t_cpx_atom_cq          (sctag0_cpx_atom_cq          ),
  .l2t_cpx_data_ca          (sctag0_cpx_data_ca[ 145 : 0 ]),
  .l2t_pcx_stall_pq         (sctag0_pcx_stall_pq         ),
  .pcx_l2t_data_rdy_px1     (pcx_sctag0_data_rdy_px1     ),
  .pcx_l2t_data_px2         (pcx_sctag0_data_px2[ 129 : 0 ]),
  .pcx_l2t_atm_px1          (pcx_sctag0_atm_px1          ),
  .cpx_l2t_grant_cx         (cpx_sctag0_grant_cx[ 7 : 0 ]    ),
  .l2t_rst_fatal_error      (l2t0_rst_fatal_error        ),
  .rst_wmr_protect                (rst_wmr_protect                 ),
  .l2t_l2d_way_sel_c2       (l2t0_l2d0_way_sel_c2        ),
  .l2t_l2d_rd_wr_c2         (l2t0_l2d0_rd_wr_c2          ),
  .l2t_l2d_set_c2           (l2t0_l2d0_set_c2[ 8 : 0 ]       ),
  .l2t_l2d_col_offset_c2    (l2t0_l2d0_col_offset_c2[ 3 : 0 ]),
  .l2t_l2d_word_en_c2       (l2t0_l2d0_word_en_c2        ),
  .l2t_l2d_fbrd_c3          (l2t0_l2d0_fbrd_c3           ),
  .l2t_l2d_fb_hit_c3        (l2t0_l2d0_fb_hit_c3         ),
  .l2t_l2d_stdecc_c2        (l2t0_l2d0_stdecc_c2[ 77 : 0 ]         ),
  .l2d_l2t_decc_c6          (l2d0_l2t0_decc_c6           ),
//  .l2t_l2b_stdecc_c3        (l2t0_l2b0_stdecc_c3[77:0]   ),
  .l2t_l2b_fbrd_en_c3       (l2t0_l2b0_fbrd_en_c3        ),
  .l2t_l2b_fbrd_wl_c3       (l2t0_l2b0_fbrd_wl_c3[ 2 : 0 ]   ),
  .l2t_l2b_fbwr_wen_r2      (l2t0_l2b0_fbwr_wen_r2[ 15 : 0 ] ),
  .l2t_l2b_fbwr_wl_r2       (l2t0_l2b0_fbwr_wl_r2[ 2 : 0 ]   ),
  .l2t_l2b_fbd_stdatasel_c3 (l2t0_l2b0_fbd_stdatasel_c3  ),
  .l2t_l2b_wbwr_wen_c6      (l2t0_l2b0_wbwr_wen_c6[ 3 : 0 ]  ),
  .l2t_l2b_wbwr_wl_c6       (l2t0_l2b0_wbwr_wl_c6[ 2 : 0 ]   ),
  .l2t_l2b_wbrd_en_r0       (l2t0_l2b0_wbrd_en_r0        ),
  .l2t_l2b_wbrd_wl_r0       (l2t0_l2b0_wbrd_wl_r0[ 2 : 0 ]   ),
  .l2t_l2b_ev_dword_r0      (l2t0_l2b0_ev_dword_r0[ 2 : 0 ]  ),
  .l2t_l2b_evict_en_r0      (l2t0_l2b0_evict_en_r0       ),
  .l2b_l2t_ev_uerr_r5       (l2b0_l2t0_ev_uerr_r5        ),
  .l2b_l2t_ev_cerr_r5       (l2b0_l2t0_ev_cerr_r5        ),
  .l2t_l2b_rdma_wren_s2     (l2t0_l2b0_rdma_wren_s2[ 15 : 0 ]),
  .l2t_l2b_rdma_wrwl_s2     (l2t0_l2b0_rdma_wrwl_s2[ 1 : 0 ] ),
  .l2t_l2b_rdma_rdwl_r0     (l2t0_l2b0_rdma_rdwl_r0[ 1 : 0 ] ),
  .l2t_l2b_rdma_rden_r0     (l2t0_l2b0_rdma_rden_r0      ),
  .l2t_l2b_ctag_en_c7       (l2t0_l2b0_ctag_en_c7        ),
  .l2t_l2b_ctag_c7          (l2t0_l2b0_ctag_c7[ 31 : 0 ]     ),
  .l2t_l2b_word_c7          (l2t0_l2b0_word_c7[ 3 : 0 ]      ),
  .l2t_l2b_req_en_c7        (l2t0_l2b0_req_en_c7         ),
  .l2t_l2b_word_vld_c7      (l2t0_l2b0_word_vld_c7       ),
  .l2b_l2t_rdma_uerr_c10    (l2b0_l2t0_rdma_uerr_c10     ),
  .l2b_l2t_rdma_cerr_c10    (l2b0_l2t0_rdma_cerr_c10     ),
  .l2b_l2t_rdma_notdata_c10 (l2b0_l2t0_rdma_notdata_c10  ),
  .l2t_mcu_rd_req           (l2t0_mcu0_rd_req            ),
  .l2t_mcu_rd_dummy_req     (l2t0_mcu0_rd_dummy_req      ),
  .l2t_mcu_rd_req_id        (l2t0_mcu0_rd_req_id[ 2 : 0 ]    ),
  .l2t_mcu_addr             (l2t0_mcu0_addr[ 39 : 7 ]        ),
  .l2t_mcu_addr_5           (l2t0_mcu0_addr_5            ),
  .l2t_mcu_wr_req           (l2t0_mcu0_wr_req            ),
  .mcu_l2t_rd_ack           (mcu0_l2t0_rd_ack            ),
  .mcu_l2t_wr_ack           (mcu0_l2t0_wr_ack            ),
  .mcu_l2t_chunk_id_r0      (mcu0_l2t0_qword_id_r0[ 1 : 0 ]  ),
  .mcu_l2t_data_vld_r0      (mcu0_l2t0_data_vld_r0       ),
  .mcu_l2t_rd_req_id_r0     (mcu0_l2t0_rd_req_id_r0[ 2 : 0 ] ),
  .mcu_l2t_secc_err_r2      (mcu0_l2t0_secc_err_r2       ),
  .mcu_l2t_mecc_err_r2      (mcu0_l2t0_mecc_err_r2       ),
  .mcu_l2t_scb_mecc_err     (mcu0_l2t0_scb_mecc_err      ),
  .mcu_l2t_scb_secc_err     (mcu0_l2t0_scb_secc_err      ),
  .sii_l2t_req_vld          (sii_l2t0_req_vld            ),
  .sii_l2t_req              (sii_l2t0_req[ 31 : 0 ]          ),
  .sii_l2b_ecc              (sii_l2b0_ecc[ 6 : 0 ]           ),
  .l2t_sii_iq_dequeue       (l2t0_sii_iq_dequeue         ),
  .l2t_sii_wib_dequeue      (l2t0_sii_wib_dequeue        ),
  .rst_por_                 ( gl_l2_por_c3t ), 
  .rst_wmr_                 ( gl_l2_wmr_c3t ), 
  .scan_in                  (tcu_soc0_scan_out           ),
  .scan_out                 (l2t0_scan_out               ),
  .efu_l2t_fuse_clr          (efu_l2t0_fuse_clr          ),                       
  .efu_l2t_fuse_xfer_en      (efu_l2t0_fuse_xfer_en      ),                       
  .efu_l2t_fuse_data         (efu_l2t0246_fuse_data      ),                       
  .l2t_efu_fuse_data         (l2t0_efu_fuse_data         ),                       
  .l2t_efu_fuse_xfer_en      (l2t0_efu_fuse_xfer_en      ),                       
  .tcu_mbist_bisi_en              (tcu_mbist_bisi_en),
  .tcu_l2t_mbist_start            (tcu_l2t0_mbist_start_t1lff),
  .tcu_l2t_mbist_scan_in          (tcu_l2t0_mbist_scan_in),
  .l2t_tcu_mbist_done             (l2t0_tcu_mbist_done),
  .l2t_tcu_mbist_fail             (l2t0_tcu_mbist_fail),
  .l2t_tcu_mbist_scan_out         (l2t0_tcu_mbist_scan_out),
  .gclk                      	  ( cmp_gclk_c3_l2t0 ), // cmp_gclk_c1_r[2]            ), 
  .tcu_clk_stop ( gl_l2t0_clk_stop ),	// staged clk_stop
  .tcu_l2t_shscan_scan_in         (tcu_l2t0_shscan_scan_in ),
  .tcu_l2t_shscan_aclk            (tcu_l2t_shscan_aclk    ),
  .tcu_l2t_shscan_bclk            (tcu_l2t_shscan_bclk    ),
  .tcu_l2t_shscan_scan_en         (tcu_l2t_shscan_scan_en ),
  .tcu_l2t_shscan_pce_ov          (tcu_l2t_shscan_pce_ov  ),
  .l2t_tcu_shscan_scan_out        (l2t0_tcu_shscan_scan_out),
  .tcu_l2t_shscan_clk_stop        (tcu_l2t0_shscan_clk_stop),
  .vnw_ary                            (L2T_VNW[ 0 ]),
  .l2t_rep_in0                        (24'b0),
  .l2t_rep_in1                        (24'b0),
  .l2t_rep_in2                        (24'b0),
  .l2t_rep_in3                        (24'b0),
  .l2t_rep_in4                        (24'b0),
  .l2t_rep_in5                        (24'b0),
  .l2t_rep_in6                        (24'b0),
  .l2t_rep_in7                        (24'b0),
  .l2t_rep_in8                        (24'b0),
  .l2t_rep_in9                        (24'b0),
  .l2t_rep_in10                       (24'b0),
  .l2t_rep_in11                       (24'b0),
  .l2t_rep_in12                       (24'b0),
  .l2t_rep_in13                       (24'b0),
  .l2t_rep_in14                       (24'b0),
  .l2t_rep_in15                       (24'b0),
  .l2t_rep_in16                       (24'b0),
  .l2t_rep_in17                       (24'b0),
  .l2t_rep_in18                       (24'b0),
  .l2t_rep_in19                       (24'b0),
  .l2t_rep_out0                       (l2t0_rep_out0_unused[ 23 : 0 ]),
  .l2t_rep_out1                       (l2t0_rep_out1_unused[ 23 : 0 ]),
  .l2t_rep_out2                       (l2t0_rep_out2_unused[ 23 : 0 ]),
  .l2t_rep_out3                       (l2t0_rep_out3_unused[ 23 : 0 ]),
  .l2t_rep_out4                       (l2t0_rep_out4_unused[ 23 : 0 ]),
  .l2t_rep_out5                       (l2t0_rep_out5_unused[ 23 : 0 ]),
  .l2t_rep_out6                       (l2t0_rep_out6_unused[ 23 : 0 ]),
  .l2t_rep_out7                       (l2t0_rep_out7_unused[ 23 : 0 ]),
  .l2t_rep_out8                       (l2t0_rep_out8_unused[ 23 : 0 ]),
  .l2t_rep_out9                       (l2t0_rep_out9_unused[ 23 : 0 ]),
  .l2t_rep_out10                      (l2t0_rep_out10_unused[ 23 : 0 ]),
  .l2t_rep_out11                      (l2t0_rep_out11_unused[ 23 : 0 ]),
  .l2t_rep_out12                      (l2t0_rep_out12_unused[ 23 : 0 ]),
  .l2t_rep_out13                      (l2t0_rep_out13_unused[ 23 : 0 ]),
  .l2t_rep_out14                      (l2t0_rep_out14_unused[ 23 : 0 ]),
  .l2t_rep_out15                      (l2t0_rep_out15_unused[ 23 : 0 ]),
  .l2t_rep_out16                      (l2t0_rep_out16_unused[ 23 : 0 ]),
  .l2t_rep_out17                      (l2t0_rep_out17_unused[ 23 : 0 ]),
  .l2t_rep_out18                      (l2t0_rep_out18_unused[ 23 : 0 ]),
  .l2t_rep_out19                      (l2t0_rep_out19_unused[ 23 : 0 ]),
  .ncu_l2t_pm(ncu_l2t_pm),
  .ncu_l2t_ba01(ncu_l2t_ba01),
  .ncu_l2t_ba23(ncu_l2t_ba23),
  .ncu_l2t_ba45(ncu_l2t_ba45),
  .ncu_l2t_ba67(ncu_l2t_ba67),
  .ncu_spc0_core_enable_status(ncu_spc0_core_enable_status),
  .ncu_spc1_core_enable_status(ncu_spc1_core_enable_status),
  .ncu_spc2_core_enable_status(ncu_spc2_core_enable_status),
  .ncu_spc3_core_enable_status(ncu_spc3_core_enable_status),
  .ncu_spc4_core_enable_status(ncu_spc4_core_enable_status),
  .ncu_spc5_core_enable_status(ncu_spc5_core_enable_status),
  .ncu_spc6_core_enable_status(ncu_spc6_core_enable_status),
  .ncu_spc7_core_enable_status(ncu_spc7_core_enable_status),
  .tcu_pce_ov(tcu_pce_ov),
  .tcu_aclk(tcu_aclk),
  .tcu_bclk(tcu_bclk),
  .tcu_scan_en(tcu_scan_en),
  .tcu_muxtest(tcu_muxtest),
  .tcu_dectest(tcu_dectest),
  .tcu_atpg_mode(tcu_atpg_mode),
  .tcu_se_scancollar_in(tcu_se_scancollar_in),
  .tcu_se_scancollar_out(tcu_se_scancollar_out),
  .tcu_array_wr_inhibit(tcu_array_wr_inhibit),
  .tcu_array_bypass(tcu_array_bypass),
  .cluster_arst_l(cluster_arst_l),
  .tcu_mbist_user_mode(tcu_mbist_user_mode)
        );
//________________________________________________________________


l2b l2b0(
  .ccu_slow_cmp_sync_en ( gl_io_cmp_sync_en_c3t0 ), // ( gl_io_cmp_sync_en_c3t ), - for int6.1
  .ccu_cmp_slow_sync_en ( gl_cmp_io_sync_en_c3t0 ), // ( gl_cmp_io_sync_en_c3t ), - for int6.1
  .select_delay_mcu ( 1'b0 ),

  .gclk                     ( cmp_gclk_c3_l2b0 ), // cmp_gclk_c0_r[1]), 
  .tcu_clk_stop ( gl_l2b0_clk_stop ),	// staged clk_stop
  .rst_por_                 (gl_l2_por_c3t0 			), // ( gl_l2_por_c3t ), - for int6.1
  .rst_wmr_                 (gl_l2_wmr_c3t0 			), // ( gl_l2_wmr_c3t ), - for int6.1
  .l2t_l2b_fbrd_en_c3       (l2t0_l2b0_fbrd_en_c3        ),// scbuf
  .l2t_l2b_fbrd_wl_c3       (l2t0_l2b0_fbrd_wl_c3        ),
  .l2t_l2b_fbwr_wen_r2      (l2t0_l2b0_fbwr_wen_r2       ),
  .l2t_l2b_fbwr_wl_r2       (l2t0_l2b0_fbwr_wl_r2        ),
  .l2t_l2b_fbd_stdatasel_c3 (l2t0_l2b0_fbd_stdatasel_c3  ),
  .l2t_l2b_stdecc_c2        (l2t0_l2d0_stdecc_c2[ 77 : 0 ]         ),
  .l2t_l2b_evict_en_r0      (l2t0_l2b0_evict_en_r0       ),
  .l2t_l2b_wbwr_wen_c6      (l2t0_l2b0_wbwr_wen_c6       ),
  .l2t_l2b_wbwr_wl_c6       (l2t0_l2b0_wbwr_wl_c6        ),
  .l2t_l2b_wbrd_en_r0       (l2t0_l2b0_wbrd_en_r0        ),
  .l2t_l2b_wbrd_wl_r0       (l2t0_l2b0_wbrd_wl_r0        ),
  .l2t_l2b_ev_dword_r0      (l2t0_l2b0_ev_dword_r0       ),
  .l2t_l2b_rdma_wren_s2     (l2t0_l2b0_rdma_wren_s2      ),
  .l2t_l2b_rdma_wrwl_s2     (l2t0_l2b0_rdma_wrwl_s2      ),
  .l2t_l2b_rdma_rden_r0     (l2t0_l2b0_rdma_rden_r0      ),
  .l2t_l2b_rdma_rdwl_r0     (l2t0_l2b0_rdma_rdwl_r0      ),
  .l2t_l2b_ctag_en_c7       (l2t0_l2b0_ctag_en_c7        ),
  .l2t_l2b_ctag_c7          (l2t0_l2b0_ctag_c7[ 31 : 0 ]     ),
  .l2t_l2b_req_en_c7        (l2t0_l2b0_req_en_c7         ),
  .l2t_l2b_word_c7          (l2t0_l2b0_word_c7           ),
  .l2t_l2b_word_vld_c7      (l2t0_l2b0_word_vld_c7       ),
  .sii_l2t_req              (sii_l2t0_req                ),
  .sii_l2b_ecc              (sii_l2b0_ecc[ 6 : 0 ]           ),
  .l2b_l2d_rvalue          (l2b0_l2d0_rvalue[ 9 : 0 ]),
  .l2b_l2d_rid             (l2b0_l2d0_rid[ 6 : 0 ]),      
  .l2b_l2d_wr_en           (l2b0_l2d0_wr_en),
  .l2b_l2d_fuse_clr        (l2b0_l2d0_fuse_clr),
  .l2d_l2b_fuse_read_data  (l2d0_l2b0_fuse_data[ 9 : 0 ]),
  .efu_l2b_fuse_data       (efu_l2b0246_fuse_data),
  .efu_l2b_fuse_xfer_en    (efu_l2b0_fuse_xfer_en),
  .efu_l2b_fuse_clr        (efu_l2b0_fuse_clr),
  .l2b_efu_fuse_xfer_en    (l2b0_efu_fuse_xfer_en),
  .l2b_efu_fuse_data       (l2b0_efu_fuse_data),
  .l2b_dbg_sio_ctag_vld	    (l2b0_dbg0_sio_ctag_vld	 ),
  .l2b_dbg_sio_ack_type	    (l2b0_dbg0_sio_ack_type	 ),
  .l2b_dbg_sio_ack_dest	    (l2b0_dbg0_sio_ack_dest	 ),
  .l2b_sio_ctag_vld         (l2b0_sio_ctag_vld           ),
  .l2b_sio_data             (l2b0_sio_data[ 31 : 0 ]         ),
  .l2b_sio_parity           (l2b0_sio_parity[ 1 : 0 ]        ),     
  .l2b_sio_ue_err           (l2b0_sio_ue_err             ),
  .l2b_l2t_rdma_uerr_c10    (l2b0_l2t0_rdma_uerr_c10     ),
  .l2b_l2t_rdma_cerr_c10    (l2b0_l2t0_rdma_cerr_c10     ),
  .l2b_l2t_rdma_notdata_c10 (l2b0_l2t0_rdma_notdata_c10  ),
  .l2b_l2t_ev_uerr_r5       (l2b0_l2t0_ev_uerr_r5        ),
  .l2b_l2t_ev_cerr_r5       (l2b0_l2t0_ev_cerr_r5        ),
  .l2d_l2b_decc_out_c7      (l2d0_l2b0_decc_out_c7       ),
  .l2b_l2d_fbdecc_c4        (l2b0_l2d0_fbdecc_c4         ),
  .mcu_l2b_data_r2          (mcu0_l2b01_data_r2[ 127 : 0 ]   ),
  .mcu_l2b_ecc_r2           (mcu0_l2b01_ecc_r2[ 27 : 0 ]     ),
  .tcu_mbist_bisi_en        (tcu_mbist_bisi_en           ),
  .tcu_l2b_mbist_start      (tcu_l2b0_mbist_start_ccxlff        ),
  .l2b_tcu_mbist_done       (l2b0_tcu_mbist_done         ),
  .l2b_tcu_mbist_fail       (l2b0_tcu_mbist_fail         ),
  .tcu_l2b_mbist_scan_in    (tcu_l2b0_mbist_scan_in      ),
  .l2b_tcu_mbist_scan_out   (l2b0_tcu_mbist_scan_out     ),
  .l2b_evict_l2b_mcu_data_mecc_r5
                            (l2b0_mcu0_data_mecc_r5      ),
  .evict_l2b_mcu_wr_data_r5 (l2b0_mcu0_wr_data_r5[ 63 : 0 ]  ),
  .evict_l2b_mcu_data_vld_r5(l2b0_mcu0_data_vld_r5       ),
  .scan_in                  (tcu_soch_scan_out           ),
  .scan_out                 (l2b0_scan_out               ),
  .rst_wmr_protect(rst_wmr_protect),
  .tcu_pce_ov(tcu_pce_ov),
  .tcu_aclk(tcu_aclk),
  .tcu_bclk(tcu_bclk),
  .tcu_scan_en(tcu_scan_en),
  .tcu_muxtest(tcu_muxtest),
  .tcu_dectest(tcu_dectest),
  .tcu_se_scancollar_in(tcu_se_scancollar_in),
  .tcu_se_scancollar_out(tcu_se_scancollar_out),
  .tcu_array_wr_inhibit(tcu_array_wr_inhibit),
  .tcu_atpg_mode(tcu_atpg_mode),
  .tcu_array_bypass(tcu_array_bypass),
  .cluster_arst_l(cluster_arst_l),
  .tcu_mbist_user_mode(tcu_mbist_user_mode)
//.so                       (                            )
        );
//________________________________________________________________


mcu mcu1(
  .gclk                     ( cmp_gclk_c4_mcu1 ), // cmp_gclk_c0_r[3]            ) , 
  .tcu_mcu_dr_clk_stop	( gl_mcu1_dr_clk_stop ),	// staged clk_stop
  .tcu_mcu_clk_stop	( gl_mcu1_clk_stop ),	// staged clk_stop
  .tcu_mcu_io_clk_stop	( gl_mcu1_io_clk_stop ),	// staged clk_stop
  .ccu_io_out	( gl_io_out_c3t ),	// staged div phase
  .ccu_dr_sync_en (gl_dr_sync_en_c3t),		
  .ccu_io_cmp_sync_en ( gl_io_cmp_sync_en_c3t ), 
  .ccu_cmp_io_sync_en ( gl_cmp_io_sync_en_c3t ),
  .dr_gclk                  ( dr_gclk_c4_mcu1 ), // dr_gclk_c0_r[3]             ) , 
  .tcu_mcu_fbd_clk_stop     (tcu_mcu1_fbd_clk_stop       ),
  .mcu_dbg1_rd_req_in_0	    (mcu1_dbg1_rd_req_in_0[ 3 : 0 ]  ),
  .mcu_dbg1_rd_req_in_1	    (mcu1_dbg1_rd_req_in_1[ 3 : 0 ]  ),
  .mcu_dbg1_rd_req_out	    (mcu1_dbg1_rd_req_out[ 4 : 0 ]   ),
  .mcu_dbg1_wr_req_in_0	    (mcu1_dbg1_wr_req_in_0       ),
  .mcu_dbg1_wr_req_in_1	    (mcu1_dbg1_wr_req_in_1       ),
  .mcu_dbg1_wr_req_out	    (mcu1_dbg1_wr_req_out[ 1 : 0 ]   ),
  .mcu_dbg1_mecc_err	    (mcu1_dbg1_mecc_err          ),
  .mcu_dbg1_secc_err	    (mcu1_dbg1_secc_err          ),
  .mcu_dbg1_fbd_err	    (mcu1_dbg1_fbd_err           ),
  .mcu_dbg1_err_mode	    (mcu1_dbg1_err_mode          ),
  .mcu_dbg1_err_event	    (mcu1_dbg1_err_event         ), 
  .mcu_dbg1_crc21	    (mcu1_dbg1_crc21             ),
  .l2t0_mcu_rd_req          (l2t2_mcu1_rd_req            ),
  .l2t0_mcu_wr_req          (l2t2_mcu1_wr_req            ),
  .l2t0_mcu_rd_dummy_req    (l2t2_mcu1_rd_dummy_req      ),
  .l2t0_mcu_rd_req_id       (l2t2_mcu1_rd_req_id[ 2 : 0 ]    ),
  .l2t0_mcu_addr_39to7      (l2t2_mcu1_addr[ 39 : 7 ]        ),
  .l2t0_mcu_addr_5          (l2t2_mcu1_addr_5            ),
  .mcu_l2t0_rd_ack          (mcu1_l2t2_rd_ack            ),
  .mcu_l2t0_wr_ack          (mcu1_l2t2_wr_ack            ),
  .mcu_l2t0_data_vld_r0     (mcu1_l2t2_data_vld_r0       ),
  .mcu_l2t0_rd_req_id_r0    (mcu1_l2t2_rd_req_id_r0[ 2 : 0 ] ),
  .mcu_l2t0_secc_err_r3     (mcu1_l2t2_secc_err_r2       ),
  .mcu_l2t0_mecc_err_r3     (mcu1_l2t2_mecc_err_r2       ),
  .mcu_l2t0_scb_secc_err    (mcu1_l2t2_scb_secc_err      ),
  .mcu_l2t0_scb_mecc_err    (mcu1_l2t2_scb_mecc_err      ),
  .mcu_l2t0_qword_id_r0     (mcu1_l2t2_qword_id_r0[ 1 : 0 ]  ),
  .l2t1_mcu_rd_req          (l2t3_mcu1_rd_req_t2lff            ),
  .l2t1_mcu_wr_req          (l2t3_mcu1_wr_req_t2lff            ),
  .l2t1_mcu_rd_dummy_req    (l2t3_mcu1_rd_dummy_req_t2lff      ),
  .l2t1_mcu_rd_req_id       (l2t3_mcu1_rd_req_id_t2lff[ 2 : 0 ]    ),
  .l2t1_mcu_addr_39to7      (l2t3_mcu1_addr_t2lff[ 39 : 7 ]        ),
  .l2t1_mcu_addr_5          (l2t3_mcu1_addr_5_t2lff            ),
  .mcu_l2t1_rd_ack          (mcu1_l2t3_rd_ack            ),
  .mcu_l2t1_wr_ack          (mcu1_l2t3_wr_ack            ),
  .mcu_l2t1_data_vld_r0     (mcu1_l2t3_data_vld_r0       ),
  .mcu_l2t1_rd_req_id_r0    (mcu1_l2t3_rd_req_id_r0[ 2 : 0 ] ),
  .mcu_l2t1_secc_err_r3     (mcu1_l2t3_secc_err_r2       ),
  .mcu_l2t1_mecc_err_r3     (mcu1_l2t3_mecc_err_r2       ),
  .mcu_l2t1_scb_secc_err    (mcu1_l2t3_scb_secc_err      ),
  .mcu_l2t1_scb_mecc_err    (mcu1_l2t3_scb_mecc_err      ),
  .mcu_l2t1_qword_id_r0     (mcu1_l2t3_qword_id_r0[ 1 : 0 ]  ),
  .mcu_l2b_data_r3          (mcu1_l2b23_data_r2[ 127 : 0 ]   ),
  .mcu_l2b_ecc_r3           (mcu1_l2b23_ecc_r2[ 27 : 0 ]     ),
  .l2b0_mcu_data_mecc_r5    (l2b2_mcu1_data_mecc_r5      ),
  .l2b0_mcu_wr_data_r5      (l2b2_mcu1_wr_data_r5[ 63 : 0 ]  ),
  .l2b0_mcu_data_vld_r5     (l2b2_mcu1_data_vld_r5       ),
  .l2b1_mcu_data_mecc_r5    (l2b3_mcu1_data_mecc_r5      ),
  .l2b1_mcu_wr_data_r5      (l2b3_mcu1_wr_data_r5[ 63 : 0 ]  ),
  .l2b1_mcu_data_vld_r5     (l2b3_mcu1_data_vld_r5       ),
  .mcu_pt_sync_out          (mcu1_pt_sync_out            ),
  .mcu_pt_sync_in0          (mcu2_pt_sync_out            ),
  .mcu_pt_sync_in1          (mcu3_pt_sync_out            ),
  .mcu_pt_sync_in2          (mcu0_pt_sync_out            ),
  .mcu_ncu_data             (mcu1_ncu_data[ 3 : 0 ]          ),
  .mcu_ncu_stall            (mcu1_ncu_stall              ),
  .mcu_ncu_vld              (mcu1_ncu_vld                ),
  .ncu_mcu_data             (ncu_mcu1_data[ 3 : 0 ]          ),
  .ncu_mcu_stall            (ncu_mcu1_stall              ),
  .ncu_mcu_vld              (ncu_mcu1_vld                ),
  .mcu_ncu_ecc              (mcu1_ncu_ecc                ),
  .mcu_ncu_fbr              (mcu1_ncu_fbr                ),
  .ncu_mcu_ecci             (ncu_mcu1_ecci               ),
  .ncu_mcu_fbui             (ncu_mcu1_fbui               ),
  .ncu_mcu_fbri             (ncu_mcu1_fbri               ),
  .mcu_fsr0_data            (mcu1_fsr2_data[ 119 : 0 ]       ),
  .mcu_fsr1_data            (mcu1_fsr3_data[ 119 : 0 ]       ),
  .mcu_fsr0_cfgpll_enpll    (mcu1_fsr2_cfgpll_enpll      ),
  .mcu_fsr1_cfgpll_enpll    (mcu1_fsr3_cfgpll_enpll      ),
  .mcu_fsr01_cfgpll_lb      (mcu1_fsr23_cfgpll_lb[ 1 : 0 ]   ),
  .mcu_fsr01_cfgpll_mpy     (mcu1_fsr23_cfgpll_mpy[ 3 : 0 ]  ),
  .mcu_fsr0_cfgrx_enrx      (mcu1_fsr2_cfgrx_enrx        ),
  .mcu_fsr1_cfgrx_enrx      (mcu1_fsr3_cfgrx_enrx        ),
  .mcu_fsr0_cfgrx_align     (mcu1_fsr2_cfgrx_align       ),
  .mcu_fsr1_cfgrx_align     (mcu1_fsr3_cfgrx_align       ),
  .mcu_fsr0_cfgrx_invpair   (mcu1_fsr2_cfgrx_invpair[ 13 : 0 ]),
  .mcu_fsr1_cfgrx_invpair   (mcu1_fsr3_cfgrx_invpair[ 13 : 0 ]),
  .mcu_fsr01_cfgrx_eq       (mcu1_fsr23_cfgrx_eq[ 3 : 0 ]    ),
  .mcu_fsr01_cfgrx_cdr      (mcu1_fsr23_cfgrx_cdr[ 2 : 0 ]   ),
  .mcu_fsr01_cfgrx_term     (mcu1_fsr23_cfgrx_term[ 2 : 0 ]  ),
  .mcu_fsr0_cfgtx_entx      (mcu1_fsr2_cfgtx_entx        ),
  .mcu_fsr1_cfgtx_entx      (mcu1_fsr3_cfgtx_entx        ),
  .mcu_fsr0_cfgtx_enidl     (mcu1_fsr2_cfgtx_enidl       ),
  .mcu_fsr1_cfgtx_enidl     (mcu1_fsr3_cfgtx_enidl       ),
  .mcu_fsr0_cfgtx_invpair   (mcu1_fsr2_cfgtx_invpair[ 9 : 0 ]),
  .mcu_fsr1_cfgtx_invpair   (mcu1_fsr3_cfgtx_invpair[ 9 : 0 ]),
  .mcu_fsr01_cfgtx_enftp    (mcu1_fsr23_cfgtx_enftp      ),
  .mcu_fsr01_cfgtx_de       (mcu1_fsr23_cfgtx_de[ 3 : 0 ]    ),
  .mcu_fsr01_cfgtx_swing    (mcu1_fsr23_cfgtx_swing[ 2 : 0 ] ),
  .mcu_fsr01_cfgtx_cm       (mcu1_fsr23_cfgtx_cm         ),
  .mcu_fsr01_cfgrtx_rate    (mcu1_fsr23_cfgrtx_rate[ 1 : 0 ] ),
  .mcu_fsr0_cfgrx_entest    (mcu1_fsr2_cfgrx_entest      ),
  .mcu_fsr1_cfgrx_entest    (mcu1_fsr3_cfgrx_entest      ),
  .mcu_fsr0_cfgtx_entest    (mcu1_fsr2_cfgtx_entest      ),
  .mcu_fsr1_cfgtx_entest    (mcu1_fsr3_cfgtx_entest      ),
  .mcu_fsr0_cfgtx_bstx      (mcu1_fsr2_cfgtx_bstx[ 9 : 0 ]   ),
  .mcu_fsr1_cfgtx_bstx      (mcu1_fsr3_cfgtx_bstx[ 9 : 0 ]   ),
  .fsr0_mcu_data            (fsr2_mcu1_data[ 167 : 0 ]       ),
  .fsr1_mcu_data            (fsr3_mcu1_data[ 167 : 0 ]       ),
  .fsr0_mcu_rxbclk          (fsr2_mcu1_rxbclk[ 13 : 0 ]      ),
  .fsr1_mcu_rxbclk          (fsr3_mcu1_rxbclk[ 13 : 0 ]      ),
  .fsr0_mcu_stspll_lock     (fsr2_mcu1_stspll_lock[ 2 : 0 ]  ),
  .fsr1_mcu_stspll_lock     (fsr3_mcu1_stspll_lock[ 2 : 0 ]  ),
  .mcu_fsr0_testcfg         (mcu1_fsr2_testcfg[ 11 : 0 ]     ),
  .mcu_fsr1_testcfg         (mcu1_fsr3_testcfg[ 11 : 0 ]     ),
  .fsr0_mcu_stsrx_sync      ({fsr2_mcu1_stsrx_sync[ 8 ],    fsr2_mcu1_stsrx_sync[ 9 ],
			      fsr2_mcu1_stsrx_sync[ 13 : 10 ],fsr2_mcu1_stsrx_sync[ 7 : 0 ]}),
  .fsr1_mcu_stsrx_sync      ({fsr3_mcu1_stsrx_sync[ 8 ],    fsr3_mcu1_stsrx_sync[ 9 ],
			      fsr3_mcu1_stsrx_sync[ 13 : 10 ],fsr3_mcu1_stsrx_sync[ 7 : 0 ]}),
  .fsr0_mcu_stsrx_losdtct   ({fsr2_mcu1_stsrx_losdtct[ 8 ],    fsr2_mcu1_stsrx_losdtct[ 9 ],
			      fsr2_mcu1_stsrx_losdtct[ 13 : 10 ],fsr2_mcu1_stsrx_losdtct[ 7 : 0 ]}),
  .fsr1_mcu_stsrx_losdtct   ({fsr3_mcu1_stsrx_losdtct[ 8 ],    fsr3_mcu1_stsrx_losdtct[ 9 ],
			      fsr3_mcu1_stsrx_losdtct[ 13 : 10 ],fsr3_mcu1_stsrx_losdtct[ 7 : 0 ]}),
  .fsr0_mcu_stsrx_testfail  (fsr2_mcu1_stsrx_testfail[ 13 : 0 ]),
  .fsr1_mcu_stsrx_testfail  (fsr3_mcu1_stsrx_testfail[ 13 : 0 ]),
  .fsr0_mcu_stsrx_bsrxp     (fsr2_mcu1_stsrx_bsrxp[ 13 : 0 ] ),
  .fsr1_mcu_stsrx_bsrxp     (fsr3_mcu1_stsrx_bsrxp[ 13 : 0 ] ),
  .fsr0_mcu_stsrx_bsrxn     (fsr2_mcu1_stsrx_bsrxn[ 13 : 0 ] ),
  .fsr1_mcu_stsrx_bsrxn     (fsr3_mcu1_stsrx_bsrxn[ 13 : 0 ] ),
  .fsr0_mcu_ststx_testfail  (fsr2_mcu1_ststx_testfail[ 9 : 0 ]),
  .fsr1_mcu_ststx_testfail  (fsr3_mcu1_ststx_testfail[ 9 : 0 ]),
  .mcu_id                   ({1'b0,1'b1}                 ),
  .tcu_mcu_mbist_start      (tcu_mcu1_mbist_start_t1lff        ),
  .mcu_tcu_mbist_done       (mcu1_tcu_mbist_done         ),
  .mcu_tcu_mbist_fail       (mcu1_tcu_mbist_fail         ),
  .tcu_mcu_mbist_scan_in    (tcu_mcu1_mbist_scan_in      ),
  .mcu_tcu_mbist_scan_out   (mcu1_tcu_mbist_scan_out     ),
  .mcu_sbs_scan_in          (mcu0_sbs_scan_out           ),
  .mcu_sbs_scan_out         (mcu1_sbs_scan_out           ),
  .scan_in                  (tcu_socc_scan_out           ),
  .scan_out                 (mcu1_scan_out               ),
  .ncu_mcu_pm(ncu_mcu_pm),
  .ncu_mcu_ba01(ncu_mcu_ba01),
  .ncu_mcu_ba23(ncu_mcu_ba23),
  .ncu_mcu_ba45(ncu_mcu_ba45),
  .ncu_mcu_ba67(ncu_mcu_ba67),
  .tcu_mbist_bisi_en(tcu_mbist_bisi_en),
  .tcu_mbist_user_mode(tcu_mbist_user_mode),
  .tcu_sbs_scan_en(tcu_sbs_scan_en),
  .tcu_sbs_aclk(tcu_sbs_aclk),
  .tcu_sbs_bclk(tcu_sbs_bclk),
  .tcu_sbs_clk(tcu_sbs_clk),
  .tcu_sbs_uclk(tcu_sbs_uclk),
  .rst_mcu_selfrsh(rst_mcu_selfrsh),
  .rst_wmr_protect(rst_wmr_protect),
  .tcu_aclk(tcu_aclk),
  .tcu_bclk(tcu_bclk),
  .tcu_pce_ov(tcu_pce_ov),
  .tcu_dectest(tcu_dectest),
  .tcu_muxtest(tcu_muxtest),
  .tcu_mcu_testmode(tcu_mcu_testmode),
  .tcu_scan_en(tcu_scan_en),
  .tcu_se_scancollar_in(tcu_se_scancollar_in),
  .tcu_array_wr_inhibit(tcu_array_wr_inhibit),
  .tcu_array_bypass(tcu_array_bypass),
  .tcu_atpg_mode(tcu_atpg_mode),
  .tcu_div_bypass(tcu_div_bypass),
  .ccu_serdes_dtm(ccu_serdes_dtm)
         );

/*
peu peu(

    .rst_por_                 (gl_dmu_peu_por_c3b ), 
    .rst_wmr_                 (gl_dmu_peu_wmr_c3b ), 
    .tcu_aclk               ( tcu_asic_aclk             ),
    .tcu_bclk               ( tcu_asic_bclk             ),
    .tcu_scan_en            ( tcu_asic_scan_en          ),
    .tcu_se_scancollar_in   ( tcu_asic_se_scancollar_in ),
    .tcu_array_wr_inhibit   ( tcu_asic_array_wr_inhibit ),
    .scan_in                (tcu_peu_scan_out),
    .scan_out               (peu_scan_out         ), // to be connected to tcu
    .peu_sbs_scan_in        (mcu1_sbs_scan_out ),
    .peu_sbs_scan_out       (peu_mac_sbs_input ),     	//  0324

    .gclk                   ( cmp_gclk_c3_peu ), 	// cmp_gclk_c0_r[0] ), 
    .tcu_peu_io_clk_stop    ( gl_peu_io_clk_stop ),	// staged clk_stop
    .ccu_io_out	( gl_io_out_c3b ),	// staged div phase
    .pc_clk                 (psr_peu_txbclk0 ),
  .ccu_serdes_dtm(ccu_serdes_dtm),
  .cluster_arst_l(cluster_arst_l),
  .rst_dmu_async_por_(rst_dmu_async_por_),
  .tcu_pce_ov(tcu_pce_ov),
  .tcu_peu_pc_clk_stop(tcu_peu_pc_clk_stop),
  .tcu_atpg_mode(tcu_atpg_mode),
  .tcu_div_bypass(tcu_div_bypass),
  .tcu_test_protect(tcu_test_protect),
  .tcu_peu_entestcfg(tcu_peu_entestcfg),
  .tcu_peu_testmode(tcu_peu_testmode),
  .tcu_peu_clk_ext(tcu_peu_clk_ext),
  .tcu_mbist_bisi_en(tcu_mbist_bisi_en),
  .tcu_mbist_user_mode(tcu_mbist_user_mode),
  .tcu_peu_mbist_start(tcu_peu_mbist_start),
  .peu_tcu_mbist_done(peu_tcu_mbist_done),
  .peu_tcu_mbist_fail(peu_tcu_mbist_fail),
  .tcu_peu_mbist_scan_in(tcu_peu_mbist_scan_in),
  .peu_tcu_mbist_scan_out(peu_tcu_mbist_scan_out),
  .tcu_sbs_scan_en(tcu_sbs_scan_en),
  .tcu_sbs_aclk(tcu_sbs_aclk),
  .tcu_sbs_bclk(tcu_sbs_bclk),
  .tcu_sbs_clk(tcu_sbs_clk),
  .tcu_sbs_uclk(tcu_sbs_uclk),
  .tcu_sbs_enbstx(tcu_sbs_enbstx),
  .tcu_sbs_enbsrx(tcu_sbs_enbsrx),
  .tcu_sbs_enbspt(tcu_sbs_enbspt),
  .tcu_sbs_acmode(tcu_sbs_acmode),
  .tcu_sbs_actestsignal(tcu_sbs_actestsignal),
  .peu_mio_debug_clk(peu_mio_debug_clk),
  .peu_mio_debug_bus_a(peu_mio_debug_bus_a[7:0]),
  .peu_mio_debug_bus_b(peu_mio_debug_bus_b[7:0]),
  .peu_mio_pipe_txdata(peu_mio_pipe_txdata[63:0]),
  .peu_mio_pipe_txdatak(peu_mio_pipe_txdatak[7:0]),
  .d2p_csr_ack(d2p_csr_ack),
  .d2p_csr_rcd(d2p_csr_rcd[95:0]),
  .d2p_csr_req(d2p_csr_req),
  .d2p_cto_ack(d2p_cto_ack),
  .d2p_ech_wptr(d2p_ech_wptr[5:0]),
  .d2p_edb_addr(d2p_edb_addr[7:0]),
  .d2p_edb_data(d2p_edb_data[127:0]),
  .d2p_edb_dpar(d2p_edb_dpar[3:0]),
  .d2p_edb_we(d2p_edb_we),
  .d2p_ehb_addr(d2p_ehb_addr[5:0]),
  .d2p_ehb_data(d2p_ehb_data[127:0]),
  .d2p_ehb_dpar(d2p_ehb_dpar[3:0]),
  .d2p_ehb_we(d2p_ehb_we),
  .d2p_erh_wptr(d2p_erh_wptr[5:0]),
  .d2p_ibc_nhc(d2p_ibc_nhc[7:0]),
  .d2p_ibc_pdc(d2p_ibc_pdc[11:0]),
  .d2p_ibc_phc(d2p_ibc_phc[7:0]),
  .d2p_ibc_req(d2p_ibc_req),
  .d2p_idb_addr(d2p_idb_addr[7:0]),
  .d2p_idb_rd(d2p_idb_rd),
  .d2p_ihb_addr(d2p_ihb_addr[5:0]),
  .d2p_ihb_rd(d2p_ihb_rd),
  .d2p_req_id(d2p_req_id[15:0]),
  .d2p_spare(d2p_spare[4:0]),
  .p2d_ce_int(p2d_ce_int),
  .p2d_csr_ack(p2d_csr_ack),
  .p2d_csr_rcd(p2d_csr_rcd[95:0]),
  .p2d_csr_req(p2d_csr_req),
  .p2d_cto_req(p2d_cto_req),
  .p2d_cto_tag(p2d_cto_tag[4:0]),
  .p2d_drain(p2d_drain),
  .p2d_ecd_rptr(p2d_ecd_rptr[7:0]),
  .p2d_ech_rptr(p2d_ech_rptr[5:0]),
  .p2d_erd_rptr(p2d_erd_rptr[7:0]),
  .p2d_erh_rptr(p2d_erh_rptr[5:0]),
  .p2d_ibc_ack(p2d_ibc_ack),
  .p2d_idb_data(p2d_idb_data[127:0]),
  .p2d_idb_dpar(p2d_idb_dpar[3:0]),
  .p2d_ihb_data(p2d_ihb_data[127:0]),
  .p2d_ihb_dpar(p2d_ihb_dpar[3:0]),
  .p2d_ihb_wptr(p2d_ihb_wptr[6:0]),
  .p2d_mps(p2d_mps[2:0]),
  .p2d_oe_int(p2d_oe_int),
  .p2d_spare(p2d_spare[4:0]),
  .p2d_ue_int(p2d_ue_int),
  .p2d_npwr_stall_en(p2d_npwr_stall_en),
  .psr_peu_rd_b0sds0(psr_peu_rd_b0sds0[9:0]),
  .psr_peu_rd_b1sds0(psr_peu_rd_b1sds0[9:0]),
  .psr_peu_rd_b2sds0(psr_peu_rd_b2sds0[9:0]),
  .psr_peu_rd_b3sds0(psr_peu_rd_b3sds0[9:0]),
  .psr_peu_rd_b0sds1(psr_peu_rd_b0sds1[9:0]),
  .psr_peu_rd_b1sds1(psr_peu_rd_b1sds1[9:0]),
  .psr_peu_rd_b2sds1(psr_peu_rd_b2sds1[9:0]),
  .psr_peu_rd_b3sds1(psr_peu_rd_b3sds1[9:0]),
  .psr_peu_rxbclk_b0sds0(psr_peu_rxbclk_b0sds0),
  .psr_peu_rxbclk_b1sds0(psr_peu_rxbclk_b1sds0),
  .psr_peu_rxbclk_b2sds0(psr_peu_rxbclk_b2sds0),
  .psr_peu_rxbclk_b3sds0(psr_peu_rxbclk_b3sds0),
  .psr_peu_rxbclk_b0sds1(psr_peu_rxbclk_b0sds1),
  .psr_peu_rxbclk_b1sds1(psr_peu_rxbclk_b1sds1),
  .psr_peu_rxbclk_b2sds1(psr_peu_rxbclk_b2sds1),
  .psr_peu_rxbclk_b3sds1(psr_peu_rxbclk_b3sds1),
  .psr_peu_bsrxn_b0sds0(psr_peu_bsrxn_b0sds0),
  .psr_peu_bsrxn_b1sds0(psr_peu_bsrxn_b1sds0),
  .psr_peu_bsrxn_b2sds0(psr_peu_bsrxn_b2sds0),
  .psr_peu_bsrxn_b3sds0(psr_peu_bsrxn_b3sds0),
  .psr_peu_bsrxn_b0sds1(psr_peu_bsrxn_b0sds1),
  .psr_peu_bsrxn_b1sds1(psr_peu_bsrxn_b1sds1),
  .psr_peu_bsrxn_b2sds1(psr_peu_bsrxn_b2sds1),
  .psr_peu_bsrxn_b3sds1(psr_peu_bsrxn_b3sds1),
  .psr_peu_bsrxp_b0sds0(psr_peu_bsrxp_b0sds0),
  .psr_peu_bsrxp_b1sds0(psr_peu_bsrxp_b1sds0),
  .psr_peu_bsrxp_b2sds0(psr_peu_bsrxp_b2sds0),
  .psr_peu_bsrxp_b3sds0(psr_peu_bsrxp_b3sds0),
  .psr_peu_bsrxp_b0sds1(psr_peu_bsrxp_b0sds1),
  .psr_peu_bsrxp_b1sds1(psr_peu_bsrxp_b1sds1),
  .psr_peu_bsrxp_b2sds1(psr_peu_bsrxp_b2sds1),
  .psr_peu_bsrxp_b3sds1(psr_peu_bsrxp_b3sds1),
  .psr_peu_losdtct_b0sds0(psr_peu_losdtct_b0sds0),
  .psr_peu_losdtct_b1sds0(psr_peu_losdtct_b1sds0),
  .psr_peu_losdtct_b2sds0(psr_peu_losdtct_b2sds0),
  .psr_peu_losdtct_b3sds0(psr_peu_losdtct_b3sds0),
  .psr_peu_losdtct_b0sds1(psr_peu_losdtct_b0sds1),
  .psr_peu_losdtct_b1sds1(psr_peu_losdtct_b1sds1),
  .psr_peu_losdtct_b2sds1(psr_peu_losdtct_b2sds1),
  .psr_peu_losdtct_b3sds1(psr_peu_losdtct_b3sds1),
  .psr_peu_sync_b0sds0(psr_peu_sync_b0sds0),
  .psr_peu_sync_b1sds0(psr_peu_sync_b1sds0),
  .psr_peu_sync_b2sds0(psr_peu_sync_b2sds0),
  .psr_peu_sync_b3sds0(psr_peu_sync_b3sds0),
  .psr_peu_sync_b0sds1(psr_peu_sync_b0sds1),
  .psr_peu_sync_b1sds1(psr_peu_sync_b1sds1),
  .psr_peu_sync_b2sds1(psr_peu_sync_b2sds1),
  .psr_peu_sync_b3sds1(psr_peu_sync_b3sds1),
  .psr_peu_rx_tstfail_b0sds0(psr_peu_rx_tstfail_b0sds0),
  .psr_peu_rx_tstfail_b1sds0(psr_peu_rx_tstfail_b1sds0),
  .psr_peu_rx_tstfail_b2sds0(psr_peu_rx_tstfail_b2sds0),
  .psr_peu_rx_tstfail_b3sds0(psr_peu_rx_tstfail_b3sds0),
  .psr_peu_rx_tstfail_b0sds1(psr_peu_rx_tstfail_b0sds1),
  .psr_peu_rx_tstfail_b1sds1(psr_peu_rx_tstfail_b1sds1),
  .psr_peu_rx_tstfail_b2sds1(psr_peu_rx_tstfail_b2sds1),
  .psr_peu_rx_tstfail_b3sds1(psr_peu_rx_tstfail_b3sds1),
  .psr_peu_rdtcip_b0sds0(psr_peu_rdtcip_b0sds0),
  .psr_peu_rdtcip_b1sds0(psr_peu_rdtcip_b1sds0),
  .psr_peu_rdtcip_b2sds0(psr_peu_rdtcip_b2sds0),
  .psr_peu_rdtcip_b3sds0(psr_peu_rdtcip_b3sds0),
  .psr_peu_rdtcip_b0sds1(psr_peu_rdtcip_b0sds1),
  .psr_peu_rdtcip_b1sds1(psr_peu_rdtcip_b1sds1),
  .psr_peu_rdtcip_b2sds1(psr_peu_rdtcip_b2sds1),
  .psr_peu_rdtcip_b3sds1(psr_peu_rdtcip_b3sds1),
  .psr_peu_tx_tstfail_b0sds0(psr_peu_tx_tstfail_b0sds0),
  .psr_peu_tx_tstfail_b1sds0(psr_peu_tx_tstfail_b1sds0),
  .psr_peu_tx_tstfail_b2sds0(psr_peu_tx_tstfail_b2sds0),
  .psr_peu_tx_tstfail_b3sds0(psr_peu_tx_tstfail_b3sds0),
  .psr_peu_tx_tstfail_b0sds1(psr_peu_tx_tstfail_b0sds1),
  .psr_peu_tx_tstfail_b1sds1(psr_peu_tx_tstfail_b1sds1),
  .psr_peu_tx_tstfail_b2sds1(psr_peu_tx_tstfail_b2sds1),
  .psr_peu_tx_tstfail_b3sds1(psr_peu_tx_tstfail_b3sds1),
  .psr_peu_lock_sds0(psr_peu_lock_sds0),
  .psr_peu_lock_sds1(psr_peu_lock_sds1),
  .peu_psr_td_b0sds0(peu_psr_td_b0sds0[9:0]),
  .peu_psr_td_b1sds0(peu_psr_td_b1sds0[9:0]),
  .peu_psr_td_b2sds0(peu_psr_td_b2sds0[9:0]),
  .peu_psr_td_b3sds0(peu_psr_td_b3sds0[9:0]),
  .peu_psr_td_b0sds1(peu_psr_td_b0sds1[9:0]),
  .peu_psr_td_b1sds1(peu_psr_td_b1sds1[9:0]),
  .peu_psr_td_b2sds1(peu_psr_td_b2sds1[9:0]),
  .peu_psr_td_b3sds1(peu_psr_td_b3sds1[9:0]),
  .peu_psr_invpair_b0sds0(peu_psr_invpair_b0sds0),
  .peu_psr_invpair_b1sds0(peu_psr_invpair_b1sds0),
  .peu_psr_invpair_b2sds0(peu_psr_invpair_b2sds0),
  .peu_psr_invpair_b3sds0(peu_psr_invpair_b3sds0),
  .peu_psr_invpair_b0sds1(peu_psr_invpair_b0sds1),
  .peu_psr_invpair_b1sds1(peu_psr_invpair_b1sds1),
  .peu_psr_invpair_b2sds1(peu_psr_invpair_b2sds1),
  .peu_psr_invpair_b3sds1(peu_psr_invpair_b3sds1),
  .peu_psr_rx_lane_ctl_0(peu_psr_rx_lane_ctl_0[15:0]),
  .peu_psr_rx_lane_ctl_1(peu_psr_rx_lane_ctl_1[15:0]),
  .peu_psr_rx_lane_ctl_2(peu_psr_rx_lane_ctl_2[15:0]),
  .peu_psr_rx_lane_ctl_3(peu_psr_rx_lane_ctl_3[15:0]),
  .peu_psr_rx_lane_ctl_4(peu_psr_rx_lane_ctl_4[15:0]),
  .peu_psr_rx_lane_ctl_5(peu_psr_rx_lane_ctl_5[15:0]),
  .peu_psr_rx_lane_ctl_6(peu_psr_rx_lane_ctl_6[15:0]),
  .peu_psr_rx_lane_ctl_7(peu_psr_rx_lane_ctl_7[15:0]),
  .peu_psr_rdtct_b0sds0(peu_psr_rdtct_b0sds0[1:0]),
  .peu_psr_rdtct_b1sds0(peu_psr_rdtct_b1sds0[1:0]),
  .peu_psr_rdtct_b2sds0(peu_psr_rdtct_b2sds0[1:0]),
  .peu_psr_rdtct_b3sds0(peu_psr_rdtct_b3sds0[1:0]),
  .peu_psr_rdtct_b0sds1(peu_psr_rdtct_b0sds1[1:0]),
  .peu_psr_rdtct_b1sds1(peu_psr_rdtct_b1sds1[1:0]),
  .peu_psr_rdtct_b2sds1(peu_psr_rdtct_b2sds1[1:0]),
  .peu_psr_rdtct_b3sds1(peu_psr_rdtct_b3sds1[1:0]),
  .peu_psr_enidl_b0sds0(peu_psr_enidl_b0sds0),
  .peu_psr_enidl_b1sds0(peu_psr_enidl_b1sds0),
  .peu_psr_enidl_b2sds0(peu_psr_enidl_b2sds0),
  .peu_psr_enidl_b3sds0(peu_psr_enidl_b3sds0),
  .peu_psr_enidl_b0sds1(peu_psr_enidl_b0sds1),
  .peu_psr_enidl_b1sds1(peu_psr_enidl_b1sds1),
  .peu_psr_enidl_b2sds1(peu_psr_enidl_b2sds1),
  .peu_psr_enidl_b3sds1(peu_psr_enidl_b3sds1),
  .peu_psr_bstx_b0sds0(peu_psr_bstx_b0sds0),
  .peu_psr_bstx_b1sds0(peu_psr_bstx_b1sds0),
  .peu_psr_bstx_b2sds0(peu_psr_bstx_b2sds0),
  .peu_psr_bstx_b3sds0(peu_psr_bstx_b3sds0),
  .peu_psr_bstx_b0sds1(peu_psr_bstx_b0sds1),
  .peu_psr_bstx_b1sds1(peu_psr_bstx_b1sds1),
  .peu_psr_bstx_b2sds1(peu_psr_bstx_b2sds1),
  .peu_psr_bstx_b3sds1(peu_psr_bstx_b3sds1),
  .peu_psr_tx_lane_ctl_0(peu_psr_tx_lane_ctl_0[9:0]),
  .peu_psr_tx_lane_ctl_1(peu_psr_tx_lane_ctl_1[9:0]),
  .peu_psr_tx_lane_ctl_2(peu_psr_tx_lane_ctl_2[9:0]),
  .peu_psr_tx_lane_ctl_3(peu_psr_tx_lane_ctl_3[9:0]),
  .peu_psr_tx_lane_ctl_4(peu_psr_tx_lane_ctl_4[9:0]),
  .peu_psr_tx_lane_ctl_5(peu_psr_tx_lane_ctl_5[9:0]),
  .peu_psr_tx_lane_ctl_6(peu_psr_tx_lane_ctl_6[9:0]),
  .peu_psr_tx_lane_ctl_7(peu_psr_tx_lane_ctl_7[9:0]),
  .peu_psr_txbclkin(peu_psr_txbclkin[7:0]),
  .peu_psr_testcfg_sds0(peu_psr_testcfg_sds0[15:0]),
  .peu_psr_testcfg_sds1(peu_psr_testcfg_sds1[15:0]),
  .peu_psr_pll_mpy(peu_psr_pll_mpy[3:0]),
  .peu_psr_pll_lb(peu_psr_pll_lb[1:0]) 
        );
*/
`endif
`endif  // OPENSPARC_CMP


/*
// leave this instance out of cmp model
`ifdef OPENSPARC_CMP
`else
psr psr (

   .VDDT                		(VDDT_PSR),
   .VDDD                		(VDDD_PSR),
   .VDDC                		(VDDC_PSR),
   .VDDA                		(VDDA_PSR),
   .VDDR                		(VDDR_PSR),
   .VSSA                		(VSSA_PSR),
   .dmu_psr_rate_scale_rx_b0sds0	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_rx_b1sds0	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_rx_b2sds0	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_rx_b3sds0	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_rx_b0sds1	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_rx_b1sds1	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_rx_b2sds1	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_rx_b3sds1	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_tx_b0sds0	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_tx_b1sds0	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_tx_b2sds0	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_tx_b3sds0	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_tx_b0sds1	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_tx_b1sds1	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_tx_b2sds1	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .dmu_psr_rate_scale_tx_b3sds1	(dmu_psr_rate_scale[ 1 : 0 ] ),
   .tcu_srd_atpgse_sds0			(tcu_srd_atpgse ),
   .tcu_srd_atpgmode_sds0		(tcu_srd_atpgmode[ 2 : 0 ] ),
   .tcu_srd_atpgse_sds1			(tcu_srd_atpgse ),
   .tcu_srd_atpgmode_sds1		(tcu_srd_atpgmode[ 2 : 0 ] ),
   .peu_psr_pll_mpy_sds0		(peu_psr_pll_mpy[ 3 : 0 ] ),
   .peu_psr_pll_lb_sds0			(peu_psr_pll_lb[ 1 : 0 ] ),
   .peu_psr_pll_mpy_sds1		(peu_psr_pll_mpy[ 3 : 0 ] ),
   .peu_psr_pll_lb_sds1			(peu_psr_pll_lb[ 1 : 0 ] ),
   .bsinitclk_sds0	    		(tcu_sbs_bsinitclk ) ,
   .bsinitclk_sds1	    		(tcu_sbs_bsinitclk ) ,
   .tcu_stciclk_sds0			(tcu_stciclk ),
   .tcu_stcicfg_sds0			(tcu_stcicfg[ 1 : 0 ] ),
   .tcu_stciclk_sds1			(tcu_stciclk ),
   .tcu_stcicfg_sds1			(tcu_stcicfg[ 1 : 0 ] ),
   .psr_stcid_sds0			(fsr3_stciq[ 2 ] ),
   .psr_stciq_sds0			(psr_stciq_sds0 ),
   .psr_stcid_sds1			(psr_stciq_sds0 ),
   .psr_stciq_sds1			(esr_stcid ),
   .efu_psr_fclk_sds0			(efu_psr_fclk ),
   .efu_psr_fclrz_sds0			(efu_psr_fclrz ),
   .efu_psr_fclk_sds1			(efu_psr_fclk ),
   .efu_psr_fclrz_sds1			(efu_psr_fclrz ),
   .psr_fdi_sds0			(efu_psr_fdi ),
   .psr_fdo_sds0			(psr_fdo_sds0 ),
   .psr_fdi_sds1			(psr_fdo_sds0 ),
   .psr_fdo_sds1			(psr_efu_fdo ),
   .mio_psr_testclkr_sds0		(mio_psr_testclkr ),
   .mio_psr_testclkt_sds0		(mio_psr_testclkt ),
   .mio_psr_testclkr_sds1		(mio_psr_testclkr ),
   .mio_psr_testclkt_sds1		(mio_psr_testclkt ),

// Int 6.1: Short RXBCLKIN to RXBCLK per I/O, Clk team resolution.
   .peu_psr_rxbclkin	    ({ psr_peu_rxbclk_b3sds1, psr_peu_rxbclk_b2sds1, 
			       psr_peu_rxbclk_b1sds1, psr_peu_rxbclk_b0sds1, 
			       psr_peu_rxbclk_b3sds0, psr_peu_rxbclk_b2sds0, 
			       psr_peu_rxbclk_b1sds0, psr_peu_rxbclk_b0sds0 } ),
   .psr_atpgd               		(fsr_left_atpgq ) ,         
   .psr_atpgq				(esr_atpgd ),
  .PEX_RX_N(PEX_RX_N[7:0]),
  .PEX_RX_P(PEX_RX_P[7:0]),
  .PEX_REFCLK_N(PEX_REFCLK_N),
  .PEX_REFCLK_P(PEX_REFCLK_P),
  .dmu_psr_pll_en_sds0(dmu_psr_pll_en_sds0),
  .dmu_psr_pll_en_sds1(dmu_psr_pll_en_sds1),
  .dmu_psr_rx_en_b0_sds0(dmu_psr_rx_en_b0_sds0),
  .dmu_psr_rx_en_b1_sds0(dmu_psr_rx_en_b1_sds0),
  .dmu_psr_rx_en_b2_sds0(dmu_psr_rx_en_b2_sds0),
  .dmu_psr_rx_en_b3_sds0(dmu_psr_rx_en_b3_sds0),
  .dmu_psr_rx_en_b0_sds1(dmu_psr_rx_en_b0_sds1),
  .dmu_psr_rx_en_b1_sds1(dmu_psr_rx_en_b1_sds1),
  .dmu_psr_rx_en_b2_sds1(dmu_psr_rx_en_b2_sds1),
  .dmu_psr_rx_en_b3_sds1(dmu_psr_rx_en_b3_sds1),
  .dmu_psr_tx_en_b0_sds0(dmu_psr_tx_en_b0_sds0),
  .dmu_psr_tx_en_b1_sds0(dmu_psr_tx_en_b1_sds0),
  .dmu_psr_tx_en_b2_sds0(dmu_psr_tx_en_b2_sds0),
  .dmu_psr_tx_en_b3_sds0(dmu_psr_tx_en_b3_sds0),
  .dmu_psr_tx_en_b0_sds1(dmu_psr_tx_en_b0_sds1),
  .dmu_psr_tx_en_b1_sds1(dmu_psr_tx_en_b1_sds1),
  .dmu_psr_tx_en_b2_sds1(dmu_psr_tx_en_b2_sds1),
  .dmu_psr_tx_en_b3_sds1(dmu_psr_tx_en_b3_sds1),
  .peu_psr_td_b0sds0(peu_psr_td_b0sds0[9:0]),
  .peu_psr_td_b1sds0(peu_psr_td_b1sds0[9:0]),
  .peu_psr_td_b2sds0(peu_psr_td_b2sds0[9:0]),
  .peu_psr_td_b3sds0(peu_psr_td_b3sds0[9:0]),
  .peu_psr_td_b0sds1(peu_psr_td_b0sds1[9:0]),
  .peu_psr_td_b1sds1(peu_psr_td_b1sds1[9:0]),
  .peu_psr_td_b2sds1(peu_psr_td_b2sds1[9:0]),
  .peu_psr_td_b3sds1(peu_psr_td_b3sds1[9:0]),
  .peu_psr_invpair_b0sds0(peu_psr_invpair_b0sds0),
  .peu_psr_invpair_b1sds0(peu_psr_invpair_b1sds0),
  .peu_psr_invpair_b2sds0(peu_psr_invpair_b2sds0),
  .peu_psr_invpair_b3sds0(peu_psr_invpair_b3sds0),
  .peu_psr_invpair_b0sds1(peu_psr_invpair_b0sds1),
  .peu_psr_invpair_b1sds1(peu_psr_invpair_b1sds1),
  .peu_psr_invpair_b2sds1(peu_psr_invpair_b2sds1),
  .peu_psr_invpair_b3sds1(peu_psr_invpair_b3sds1),
  .peu_psr_rx_lane_ctl_0(peu_psr_rx_lane_ctl_0[15:0]),
  .peu_psr_rx_lane_ctl_1(peu_psr_rx_lane_ctl_1[15:0]),
  .peu_psr_rx_lane_ctl_2(peu_psr_rx_lane_ctl_2[15:0]),
  .peu_psr_rx_lane_ctl_3(peu_psr_rx_lane_ctl_3[15:0]),
  .peu_psr_rx_lane_ctl_4(peu_psr_rx_lane_ctl_4[15:0]),
  .peu_psr_rx_lane_ctl_5(peu_psr_rx_lane_ctl_5[15:0]),
  .peu_psr_rx_lane_ctl_6(peu_psr_rx_lane_ctl_6[15:0]),
  .peu_psr_rx_lane_ctl_7(peu_psr_rx_lane_ctl_7[15:0]),
  .peu_psr_rdtct_b0sds0(peu_psr_rdtct_b0sds0[1:0]),
  .peu_psr_rdtct_b1sds0(peu_psr_rdtct_b1sds0[1:0]),
  .peu_psr_rdtct_b2sds0(peu_psr_rdtct_b2sds0[1:0]),
  .peu_psr_rdtct_b3sds0(peu_psr_rdtct_b3sds0[1:0]),
  .peu_psr_rdtct_b0sds1(peu_psr_rdtct_b0sds1[1:0]),
  .peu_psr_rdtct_b1sds1(peu_psr_rdtct_b1sds1[1:0]),
  .peu_psr_rdtct_b2sds1(peu_psr_rdtct_b2sds1[1:0]),
  .peu_psr_rdtct_b3sds1(peu_psr_rdtct_b3sds1[1:0]),
  .peu_psr_enidl_b0sds0(peu_psr_enidl_b0sds0),
  .peu_psr_enidl_b1sds0(peu_psr_enidl_b1sds0),
  .peu_psr_enidl_b2sds0(peu_psr_enidl_b2sds0),
  .peu_psr_enidl_b3sds0(peu_psr_enidl_b3sds0),
  .peu_psr_enidl_b0sds1(peu_psr_enidl_b0sds1),
  .peu_psr_enidl_b1sds1(peu_psr_enidl_b1sds1),
  .peu_psr_enidl_b2sds1(peu_psr_enidl_b2sds1),
  .peu_psr_enidl_b3sds1(peu_psr_enidl_b3sds1),
  .peu_psr_bstx_b0sds0(peu_psr_bstx_b0sds0),
  .peu_psr_bstx_b1sds0(peu_psr_bstx_b1sds0),
  .peu_psr_bstx_b2sds0(peu_psr_bstx_b2sds0),
  .peu_psr_bstx_b3sds0(peu_psr_bstx_b3sds0),
  .peu_psr_bstx_b0sds1(peu_psr_bstx_b0sds1),
  .peu_psr_bstx_b1sds1(peu_psr_bstx_b1sds1),
  .peu_psr_bstx_b2sds1(peu_psr_bstx_b2sds1),
  .peu_psr_bstx_b3sds1(peu_psr_bstx_b3sds1),
  .peu_psr_tx_lane_ctl_0(peu_psr_tx_lane_ctl_0[9:0]),
  .peu_psr_tx_lane_ctl_1(peu_psr_tx_lane_ctl_1[9:0]),
  .peu_psr_tx_lane_ctl_2(peu_psr_tx_lane_ctl_2[9:0]),
  .peu_psr_tx_lane_ctl_3(peu_psr_tx_lane_ctl_3[9:0]),
  .peu_psr_tx_lane_ctl_4(peu_psr_tx_lane_ctl_4[9:0]),
  .peu_psr_tx_lane_ctl_5(peu_psr_tx_lane_ctl_5[9:0]),
  .peu_psr_tx_lane_ctl_6(peu_psr_tx_lane_ctl_6[9:0]),
  .peu_psr_tx_lane_ctl_7(peu_psr_tx_lane_ctl_7[9:0]),
  .peu_psr_txbclkin(peu_psr_txbclkin[7:0]),
  .peu_psr_testcfg_sds0(peu_psr_testcfg_sds0[15:0]),
  .peu_psr_testcfg_sds1(peu_psr_testcfg_sds1[15:0]),
  .PEX_TX_N(PEX_TX_N[7:0]),
  .PEX_TX_P(PEX_TX_P[7:0]),
  .PEX_AMUX(PEX_AMUX[1:0]),
  .psr_peu_rd_b0sds0(psr_peu_rd_b0sds0[9:0]),
  .psr_peu_rd_b1sds0(psr_peu_rd_b1sds0[9:0]),
  .psr_peu_rd_b2sds0(psr_peu_rd_b2sds0[9:0]),
  .psr_peu_rd_b3sds0(psr_peu_rd_b3sds0[9:0]),
  .psr_peu_rd_b0sds1(psr_peu_rd_b0sds1[9:0]),
  .psr_peu_rd_b1sds1(psr_peu_rd_b1sds1[9:0]),
  .psr_peu_rd_b2sds1(psr_peu_rd_b2sds1[9:0]),
  .psr_peu_rd_b3sds1(psr_peu_rd_b3sds1[9:0]),
  .psr_peu_rxbclk_b0sds0(psr_peu_rxbclk_b0sds0),
  .psr_peu_rxbclk_b1sds0(psr_peu_rxbclk_b1sds0),
  .psr_peu_rxbclk_b2sds0(psr_peu_rxbclk_b2sds0),
  .psr_peu_rxbclk_b3sds0(psr_peu_rxbclk_b3sds0),
  .psr_peu_rxbclk_b0sds1(psr_peu_rxbclk_b0sds1),
  .psr_peu_rxbclk_b1sds1(psr_peu_rxbclk_b1sds1),
  .psr_peu_rxbclk_b2sds1(psr_peu_rxbclk_b2sds1),
  .psr_peu_rxbclk_b3sds1(psr_peu_rxbclk_b3sds1),
  .psr_peu_bsrxn_b0sds0(psr_peu_bsrxn_b0sds0),
  .psr_peu_bsrxn_b1sds0(psr_peu_bsrxn_b1sds0),
  .psr_peu_bsrxn_b2sds0(psr_peu_bsrxn_b2sds0),
  .psr_peu_bsrxn_b3sds0(psr_peu_bsrxn_b3sds0),
  .psr_peu_bsrxn_b0sds1(psr_peu_bsrxn_b0sds1),
  .psr_peu_bsrxn_b1sds1(psr_peu_bsrxn_b1sds1),
  .psr_peu_bsrxn_b2sds1(psr_peu_bsrxn_b2sds1),
  .psr_peu_bsrxn_b3sds1(psr_peu_bsrxn_b3sds1),
  .psr_peu_bsrxp_b0sds0(psr_peu_bsrxp_b0sds0),
  .psr_peu_bsrxp_b1sds0(psr_peu_bsrxp_b1sds0),
  .psr_peu_bsrxp_b2sds0(psr_peu_bsrxp_b2sds0),
  .psr_peu_bsrxp_b3sds0(psr_peu_bsrxp_b3sds0),
  .psr_peu_bsrxp_b0sds1(psr_peu_bsrxp_b0sds1),
  .psr_peu_bsrxp_b1sds1(psr_peu_bsrxp_b1sds1),
  .psr_peu_bsrxp_b2sds1(psr_peu_bsrxp_b2sds1),
  .psr_peu_bsrxp_b3sds1(psr_peu_bsrxp_b3sds1),
  .psr_peu_losdtct_b0sds0(psr_peu_losdtct_b0sds0),
  .psr_peu_losdtct_b1sds0(psr_peu_losdtct_b1sds0),
  .psr_peu_losdtct_b2sds0(psr_peu_losdtct_b2sds0),
  .psr_peu_losdtct_b3sds0(psr_peu_losdtct_b3sds0),
  .psr_peu_losdtct_b0sds1(psr_peu_losdtct_b0sds1),
  .psr_peu_losdtct_b1sds1(psr_peu_losdtct_b1sds1),
  .psr_peu_losdtct_b2sds1(psr_peu_losdtct_b2sds1),
  .psr_peu_losdtct_b3sds1(psr_peu_losdtct_b3sds1),
  .psr_peu_sync_b0sds0(psr_peu_sync_b0sds0),
  .psr_peu_sync_b1sds0(psr_peu_sync_b1sds0),
  .psr_peu_sync_b2sds0(psr_peu_sync_b2sds0),
  .psr_peu_sync_b3sds0(psr_peu_sync_b3sds0),
  .psr_peu_sync_b0sds1(psr_peu_sync_b0sds1),
  .psr_peu_sync_b1sds1(psr_peu_sync_b1sds1),
  .psr_peu_sync_b2sds1(psr_peu_sync_b2sds1),
  .psr_peu_sync_b3sds1(psr_peu_sync_b3sds1),
  .psr_peu_rx_tstfail_b0sds0(psr_peu_rx_tstfail_b0sds0),
  .psr_peu_rx_tstfail_b1sds0(psr_peu_rx_tstfail_b1sds0),
  .psr_peu_rx_tstfail_b2sds0(psr_peu_rx_tstfail_b2sds0),
  .psr_peu_rx_tstfail_b3sds0(psr_peu_rx_tstfail_b3sds0),
  .psr_peu_rx_tstfail_b0sds1(psr_peu_rx_tstfail_b0sds1),
  .psr_peu_rx_tstfail_b1sds1(psr_peu_rx_tstfail_b1sds1),
  .psr_peu_rx_tstfail_b2sds1(psr_peu_rx_tstfail_b2sds1),
  .psr_peu_rx_tstfail_b3sds1(psr_peu_rx_tstfail_b3sds1),
  .psr_peu_rdtcip_b0sds0(psr_peu_rdtcip_b0sds0),
  .psr_peu_rdtcip_b1sds0(psr_peu_rdtcip_b1sds0),
  .psr_peu_rdtcip_b2sds0(psr_peu_rdtcip_b2sds0),
  .psr_peu_rdtcip_b3sds0(psr_peu_rdtcip_b3sds0),
  .psr_peu_rdtcip_b0sds1(psr_peu_rdtcip_b0sds1),
  .psr_peu_rdtcip_b1sds1(psr_peu_rdtcip_b1sds1),
  .psr_peu_rdtcip_b2sds1(psr_peu_rdtcip_b2sds1),
  .psr_peu_rdtcip_b3sds1(psr_peu_rdtcip_b3sds1),
  .psr_peu_tx_tstfail_b0sds0(psr_peu_tx_tstfail_b0sds0),
  .psr_peu_tx_tstfail_b1sds0(psr_peu_tx_tstfail_b1sds0),
  .psr_peu_tx_tstfail_b2sds0(psr_peu_tx_tstfail_b2sds0),
  .psr_peu_tx_tstfail_b3sds0(psr_peu_tx_tstfail_b3sds0),
  .psr_peu_tx_tstfail_b0sds1(psr_peu_tx_tstfail_b0sds1),
  .psr_peu_tx_tstfail_b1sds1(psr_peu_tx_tstfail_b1sds1),
  .psr_peu_tx_tstfail_b2sds1(psr_peu_tx_tstfail_b2sds1),
  .psr_peu_tx_tstfail_b3sds1(psr_peu_tx_tstfail_b3sds1),
  .psr_peu_lock_sds0(psr_peu_lock_sds0),
  .psr_peu_lock_sds1(psr_peu_lock_sds1),
  .psr_peu_txbclk0(psr_peu_txbclk0) 
    );
`endif  // OPENSPARC_CMP

*/


//--------------------------------------------------------
//  added the following 5 IO modules
// // Ethernet SerDes (Called ges prior to 4-13-04.) //Replaced by real serdes

//.testcfg_a		    (24'b0			 ),
//.scancfg_a		    ( 2'b0			 ),
//.scancfg_b		    ( 2'b0			 ),
//.scanin_a		    ( 1'b0			 ),
//.testclkr_a		    ( 1'b0			 ),
//.testclkt_a		    ( 1'b0			 ),
//.bstxd_a		    ( 4'b0			 ),
//.cfg_a		    (48'b0			 ),
//.enpll_a		    ( 1'b0			 ),
//.enrx_a		    ( 4'b0			 ),
//.jogcom_a		    ( 4'b0			 ),
//.refclkn_a		    ( 1'b0			 ),
//.refclkp_a		    ( 1'b0			 ),
//.rxbclksta_a		    ( 4'b0			 ),
//.rxn0_a		    ( 1'b0			 ),
//.rxn1_a		    ( 1'b0			 ),
//.rxn2_a		    ( 1'b0			 ),
//.rxn3_a		    ( 1'b0			 ),
//.rxp0_a		    ( 1'b0			 ),
//.rxp1_a		    ( 1'b0			 ),
//.rxp2_a		    ( 1'b0			 ),
//.rxp3_a		    ( 1'b0			 ),
//.rxbclkin_a		    ( 4'b0			 ),
//.td0_a		    (10'b0			 ),
//.td1_a		    (10'b0			 ),
//.td2_a		    (10'b0			 ),
//.td3_a		    (10'b0			 ),
//.mdclk                    ( 1'b0			 ),
//.mdo                      ( 1'b0			 ),
//.mdo_0_en		    ( 1'b0			 ),
//.vref                     ( 1'b0			 ),
//.scanclk_a		    ( 1'b0			 ),
//.txbclksta_a		    ( 4'b0			 ),
//.txbclkin_a		    ( 4'b0			 ),
//.testcfg_b		    (24'b0			 ),
//.scanclk_b		    ( 1'b0			 ),
//.scanin_b		    ( 1'b0			 ),
//.testclkr_b		    ( 1'b0			 ),

//.scanin_b		    ( 1'b0			 ),
//.testclkr_b		    ( 1'b0			 ),
//.testclkt_b		    ( 1'b0			 ),
//.bstxd_b		    ( 4'b0			 ),
//.cfg_b		    (48'b0			 ),
//.enpll_b		    ( 1'b0			 ),
//.enrx_b		    ( 4'b0			 ),
//.jogcom_b		    ( 4'b0			 ),
//.refclkn_b		    ( 1'b0			 ),
//.refclkp_b		    ( 1'b0			 ),
//.rxbclksta_b		    ( 4'b0			 ),
//.rxn0_b		    ( 1'b0			 ),
//.rxn1_b		    ( 1'b0			 ),
//.rxn2_b		    ( 1'b0			 ),
//.rxn3_b		    ( 1'b0			 ),
//.rxp0_b		    ( 1'b0			 ),
//.rxp1_b		    ( 1'b0			 ),
//.rxp2_b		    ( 1'b0			 ),
//.rxp3_b		    ( 1'b0			 ),
//.rxbclkin_b		    ( 4'b0			 ),
//.td0_b		    (10'b0			 ),
//.td1_b		    (10'b0			 ),
//.td2_b		    (10'b0			 ),
//.td3_b		    (10'b0			 ),
//.txbclksta_b		    ( 4'b0			 ),
//.txbclkin_b		    ( 4'b0			 )

//	);

// leave this instance out of cmp model
`ifdef OPENSPARC_CMP
`else
rst rst (
  .scan_in                  ( tcu_rst_scan_out           ),
  .scan_out                 ( rst_scan_out               ),
//.mio_rst_pwron_rst_l      ( mio_rst_pwron_rst_l        ),// PWRON_RST_L
//.mio_rst_button_xir_l     ( mio_rst_button_xir_l       ),// BUTTON_XIR_L
//.mio_rst_pb_rst_l         ( mio_rst_pb_rst_l           ),// PB_RST_L
//.ccu_rst_sys_clk          ( ccu_rst_sys_clk            ),// Sunv name connect.
//.ccu_rst_change           ( ccu_rst_change             ),// Sunv name connect.
//.ccu_io_out               ( ccu_io_out                 ),// Sunv name connect.
  .gclk                     ( cmp_gclk_c1_db1            ), // ( cmp_gclk_c1_rst  - for int6.1 
  .ccu_io_cmp_sync_en       ( gl_io_cmp_sync_en_c1m      ), 
  .ccu_cmp_io_sync_en       ( gl_cmp_io_sync_en_c1m      ),
  .tcu_rst_io_clk_stop      ( gl_rst_io_clk_stop         ),// staged clk_stop
  .tcu_rst_clk_stop         ( gl_rst_clk_stop            ),// staged clk_stop
  .ccu_io_out               ( gl_io_out_c1m              ),
  .ccu_rst_sys_clk(ccu_rst_sys_clk),
  .tcu_div_bypass(tcu_div_bypass),
  .tcu_atpg_mode(tcu_atpg_mode),
  .tcu_pce_ov(tcu_pce_ov),
  .tcu_aclk(tcu_aclk),
  .tcu_bclk(tcu_bclk),
  .tcu_scan_en(tcu_scan_en),
  .ccu_cmp_sys_sync_en(ccu_cmp_sys_sync_en),
  .ccu_sys_cmp_sync_en(ccu_sys_cmp_sync_en),
  .ncu_rst_vld(ncu_rst_vld),
  .ncu_rst_data(ncu_rst_data[3:0]),
  .rst_ncu_stall(rst_ncu_stall),
  .rst_ncu_vld(rst_ncu_vld),
  .rst_ncu_data(rst_ncu_data[3:0]),
  .ncu_rst_stall(ncu_rst_stall),
  .mio_rst_pwron_rst_l(mio_rst_pwron_rst_l),
  .mio_rst_button_xir_l(mio_rst_button_xir_l),
  .ncu_rst_xir_done(ncu_rst_xir_done),
  .tcu_rst_flush_init_ack(tcu_rst_flush_init_ack),
  .tcu_rst_flush_stop_ack(tcu_rst_flush_stop_ack),
  .tcu_rst_asicflush_stop_ack(tcu_rst_asicflush_stop_ack),
  .mio_rst_pb_rst_l(mio_rst_pb_rst_l),
  .ccu_rst_change(ccu_rst_change),
  .tcu_bisx_done(tcu_bisx_done),
  .tcu_rst_efu_done(tcu_rst_efu_done),
  .l2t0_rst_fatal_error(l2t0_rst_fatal_error),
  .l2t1_rst_fatal_error(l2t1_rst_fatal_error),
  .l2t2_rst_fatal_error(l2t2_rst_fatal_error),
  .l2t3_rst_fatal_error(l2t3_rst_fatal_error),
  .l2t4_rst_fatal_error(l2t4_rst_fatal_error),
  .l2t5_rst_fatal_error(l2t5_rst_fatal_error),
  .l2t6_rst_fatal_error(l2t6_rst_fatal_error),
  .l2t7_rst_fatal_error(l2t7_rst_fatal_error),
  .ncu_rst_fatal_error(ncu_rst_fatal_error),
  .tcu_rst_scan_mode(tcu_rst_scan_mode),
  .ccu_rst_sync_stable(ccu_rst_sync_stable),
  .tcu_test_protect(tcu_test_protect),
  .rst_l2_por_(rst_l2_por_),
  .rst_l2_wmr_(rst_l2_wmr_),
  .rst_ccu_pll_(rst_ccu_pll_),
  .rst_ccu_(rst_ccu_),
  .rst_wmr_protect(rst_wmr_protect),
  .rst_tcu_clk_stop(rst_tcu_clk_stop),
  .rst_mcu_selfrsh(rst_mcu_selfrsh),
  .rst_tcu_flush_init_req(rst_tcu_flush_init_req),
  .rst_tcu_flush_stop_req(rst_tcu_flush_stop_req),
  .rst_tcu_asicflush_stop_req(rst_tcu_asicflush_stop_req),
  .rst_niu_mac_(rst_niu_mac_),
  .rst_niu_wmr_(rst_niu_wmr_),
  .rst_dmu_peu_por_(rst_dmu_peu_por_),
  .rst_dmu_peu_wmr_(rst_dmu_peu_wmr_),
  .rst_ncu_unpark_thread(rst_ncu_unpark_thread),
  .rst_ncu_xir_(rst_ncu_xir_),
  .rst_mio_pex_reset_l(rst_mio_pex_reset_l),
  .rst_mio_ssi_sync_l(rst_mio_ssi_sync_l),
  .rst_mio_rst_state(rst_mio_rst_state[5:0]),
  .cluster_arst_l(cluster_arst_l),
  .rst_tcu_dbr_gen(rst_tcu_dbr_gen),
  .rst_dmu_async_por_(rst_dmu_async_por_),
  .rst_tcu_pwron_rst_l(rst_tcu_pwron_rst_l)// staged div phase
        );
`endif  // OPENSPARC_CMP
//________________________________________________________________


n2_revid_cust n2_revid_cust (
   .jtag_revid_in ( 4'h3 ),
   .mask_minor    ( 4'h1 ),
  .jtag_revid_out(jtag_revid_out[3:0]),
  .spc_revid_out(spc_revid_out[3:0]));

//________________________________________________________________

n2_clk_gl_cust n2_clk_gl_cust (
	// PRIMARY INPUTS (FROM CCU) 
	.pll_dr_clk ( drl2clk ) , // .dr_pll_clk ( drl2clk ) , - for int6.1
	.pll_cmp_clk ( l2clk ) , // .cmp_pll_clk ( l2clk ) , - for int6.1
	// OTHERS -- AUTOMATIC CONNECTIONS
	// PRIMARY INPUTS (FROM RST) -- AUTOMATIC CONNECTIONS
	// PRIMARY INPUTS (FROM TCU) -- AUTOMATIC CONNECTIONS
	// STAGED INPUTS 
	.stg1_ccx_clk_stop_in_c1b ( stg1_ccx_clk_stop_c1b  ),
	.stg1_cmp_io_sync_en_in_c1b ( stg1_cmp_io_sync_en_c1b  ),
	.stg1_cmp_io_sync_en_in_c1t ( stg1_cmp_io_sync_en_c1t  ),
	.stg1_db0_clk_stop_in_c1b ( stg1_db0_clk_stop_c1b  ),
	.stg1_dmu_io_clk_stop_in_c1b ( stg1_dmu_io_clk_stop_c1b  ),
	.stg1_dmu_peu_por_in_c1b ( stg1_dmu_peu_por_c1b  ),
	.stg1_dmu_peu_wmr_in_c1b ( stg1_dmu_peu_wmr_c1b  ),
	.stg1_dr_sync_en_in_c1t ( stg1_dr_sync_en_c1t  ),
	.stg1_io2x_out_in_c1b ( stg1_io2x_out_c1b  ),
	.stg1_io_cmp_sync_en_in_c1b ( stg1_io_cmp_sync_en_c1b  ),
	.stg1_io_cmp_sync_en_in_c1t ( stg1_io_cmp_sync_en_c1t  ),
	.stg1_io_out_in_c1b ( stg1_io_out_c1b  ),
	.stg1_io_out_in_c1t ( stg1_io_out_c1t  ),
	.stg1_l2_por_in_c1b ( stg1_rst_l2_por_c1b  ),// UNDRIVEN stg1_l2_por_c1b  
	.stg1_l2_por_in_c1t ( stg1_rst_l2_por_c1t  ),// UNDRIVEN stg1_l2_por_c1t  
	.stg1_l2_wmr_in_c1b ( stg1_rst_l2_wmr_c1b  ),// UNDRIVEN stg1_l2_wmr_c1b 
	.stg1_l2_wmr_in_c1t ( stg1_rst_l2_wmr_c1t  ),// UNDRIVEN stg1_l2_wmr_c1t 
	.stg1_l2b0_clk_stop_in_c1t ( stg1_l2b0_clk_stop_c1t  ),
	.stg1_l2b1_clk_stop_in_c1t ( stg1_l2b1_clk_stop_c1t  ),
	.stg1_l2b2_clk_stop_in_c1b ( stg1_l2b2_clk_stop_c1b  ),
	.stg1_l2b3_clk_stop_in_c1b ( stg1_l2b3_clk_stop_c1b  ),
	.stg1_l2b4_clk_stop_in_c1t ( stg1_l2b4_clk_stop_c1t  ),
	.stg1_l2b5_clk_stop_in_c1t ( stg1_l2b5_clk_stop_c1t  ),
	.stg1_l2d0_clk_stop_in_c1t ( stg1_l2d0_clk_stop_c1t  ),
	.stg1_l2d1_clk_stop_in_c1t ( stg1_l2d1_clk_stop_c1t  ),
	.stg1_l2d2_clk_stop_in_c1b ( stg1_l2d2_clk_stop_c1b  ),
	.stg1_l2d3_clk_stop_in_c1b ( stg1_l2d3_clk_stop_c1b  ),
	.stg1_l2d4_clk_stop_in_c1t ( stg1_l2d4_clk_stop_c1t  ),
	.stg1_l2d5_clk_stop_in_c1t ( stg1_l2d5_clk_stop_c1t  ),
//	.stg1_l2d6_clk_stop_in_c1b ( stg1_l2d6_clk_stop_c1b  ),	// ECO1.2 	-mh157021 
	.stg1_l2d7_clk_stop_in_c1b ( stg1_l2d7_clk_stop_c1b  ), // ECO1.2	-mh157021	
	.stg1_l2t0_clk_stop_in_c1t ( stg1_l2t0_clk_stop_c1t  ),
	.stg1_l2t1_clk_stop_in_c1t ( stg1_l2t1_clk_stop_c1t  ),
	.stg1_l2t2_clk_stop_in_c1b ( stg1_l2t2_clk_stop_c1b  ),
	.stg1_l2t3_clk_stop_in_c1b ( stg1_l2t3_clk_stop_c1b  ),
	.stg1_l2t5_clk_stop_in_c1t ( stg1_l2t5_clk_stop_c1t  ),
	.stg1_l2t7_clk_stop_in_c1b ( stg1_l2t7_clk_stop_c1b  ),
	.stg1_mac_io_clk_stop_in_c1b ( stg1_mac_io_clk_stop_c1b ), // UNDRIVEN stg1_mac_clk_stop_c1b  
	.stg1_mcu0_clk_stop_in_c1t ( stg1_mcu0_clk_stop_c1t  ),
	.stg1_mcu0_dr_clk_stop_in_c2b ( stg1_mcu0_dr_clk_stop_c1t  ), // UNDRIVEN stg1_mcu0_dr_clk_stop_c2t 
	.stg1_mcu0_io_clk_stop_in_c1t ( stg1_mcu0_io_clk_stop_c1t  ),
	.stg1_mcu1_clk_stop_in_c1t ( stg1_mcu1_clk_stop_c1t  ),
	.stg1_mcu1_dr_clk_stop_in_c2b ( stg1_mcu1_dr_clk_stop_c1t  ), // UNDRIVEN stg1_mcu1_dr_clk_stop_c2t 
	.stg1_mcu1_io_clk_stop_in_c1t ( stg1_mcu1_io_clk_stop_c1t  ),
	.stg1_mio_clk_stop_in_c1t ( stg1_mio_clk_stop_c1t  ),
	.stg1_mio_io2x_sync_en_in_c1t ( stg1_io2x_sync_en_c1t ), // UNDRIVEN stg1_mio_io2x_sync_en_c1t  
	.stg1_ncu_clk_stop_in_c1b ( stg1_ncu_clk_stop_c1b  ),
	.stg1_ncu_io_clk_stop_in_c1b ( stg1_ncu_io_clk_stop_c1b  ),
	.stg1_peu_io_clk_stop_in_c1b ( stg1_peu_io_clk_stop_c1b  ),
	.stg1_rdp_io_clk_stop_in_c1b ( stg1_rdp_io_clk_stop_c1b  ), // UNDRIVEN stg1_rdp_clk_stop_c1b  
	.stg1_rst_mac_in_c1b ( stg1_rst_niu_mac_c1b ), // UNDRIVEN stg1_rst_mac_c1b  
	.stg1_rst_niu_wmr_in_c1b ( stg1_rst_niu_wmr_c1b  ),
	.stg1_tds_io_clk_stop_in_c1b (stg1_tds_io_clk_stop_c1b ), // UNDRIVEN stg1_tds_io_clk_stop_c1b  
	.stg1_rtx_io_clk_stop_in_c1b ( stg1_rtx_io_clk_stop_c1b ), // UNDRIVEN stg1_rtx_clk_stop_c1b  
	.stg1_sii_clk_stop_in_c1b ( stg1_sii_clk_stop_c1b  ),
	.stg1_sii_io_clk_stop_in_c1b ( stg1_sii_io_clk_stop_c1b  ),

	.stg1_cmp_io_sync_en_in_c1bg ( stg1_cmp_io_sync_en_c1b ), // for int6.1 (set 3)
	.stg1_cmp_io_sync_en_in_c1tg ( stg1_cmp_io_sync_en_c1t ), // for int6.1 (set 3)
	.stg1_io_cmp_sync_en_in_c1bg ( stg1_io_cmp_sync_en_c1b ), // for int6.1 (set 3)
	.stg1_io_cmp_sync_en_in_c1tg ( stg1_io_cmp_sync_en_c1t ), // for int6.1 (set 3)
	.stg1_io_out_in_c1bg ( stg1_io_out_c1b ), // for int6.1 (set 3)
	.stg1_l2_por_in_c1bg ( stg1_rst_l2_por_c1b ), // for int6.1 (set 3)
	.stg1_l2_por_in_c1tg ( stg1_rst_l2_por_c1t ), // for int6.1 (set 3)
	.stg1_l2_wmr_in_c1bg ( stg1_rst_l2_wmr_c1b ), // for int6.1 (set 3)
	.stg1_l2_wmr_in_c1tg ( stg1_rst_l2_wmr_c1t ), // for int6.1 (set 3)
	.stg1_mio_clk_stop_in_c1tg ( stg1_mio_clk_stop_c1t ), // for int6.1 (set 3)
	.stg1_mio_io2x_sync_en_in_c1tg ( stg1_io2x_sync_en_c1t ), // for int6.1 (set 3)
	.stg4_cmp_io_sync_en_in_c3t0 ( stg4_cmp_io_sync_en_c3t ), // for int6.1 (set 3)
	.stg4_io_cmp_sync_en_in_c3t0 ( stg4_io_cmp_sync_en_c3t ), // for int6.1 (set 3)
	.stg4_io_out_in_c3b0 ( stg4_io_out_c3b ), // for int6.1 (set 3)
	.stg4_l2_por_in_c3t0 ( stg4_l2_por_c3t ), // for int6.1 (set 3)
	.stg4_l2_wmr_in_c3t0 ( stg4_l2_wmr_c3t ), // for int6.1 (set 3)

	.stg1_spc0_clk_stop_in_c1t ( stg1_spc0_clk_stop_c1t  ),
	.stg1_spc1_clk_stop_in_c1t ( stg1_spc1_clk_stop_c1t  ),
	.stg1_spc2_clk_stop_in_c1b ( stg1_spc2_clk_stop_c1b  ),
	.stg1_spc3_clk_stop_in_c1b ( stg1_spc3_clk_stop_c1b  ),
	.stg1_spc4_clk_stop_in_c1t ( stg1_spc4_clk_stop_c1t  ),
	.stg1_spc5_clk_stop_in_c1t ( stg1_spc5_clk_stop_c1t  ),
	.stg1_spc6_clk_stop_in_c1b ( stg1_spc6_clk_stop_c1b  ), // for int6.1 (set 3)
	.stg1_spc7_clk_stop_in_c1b ( stg1_spc7_clk_stop_c1b  ),
	.stg2_ccx_clk_stop_in_c2b ( stg2_ccx_clk_stop_c1b  ),// UNDRIVEN stg2_ccx_clk_stop_c2b  
	.stg2_cmp_io_sync_en_in_c2b ( stg2_cmp_io_sync_en_c1b  ),// UNDRIVEN stg2_cmp_io_sync_en_c2b  
	.stg2_cmp_io_sync_en_in_c2t ( stg2_cmp_io_sync_en_c1t  ),// UNDRIVEN stg2_cmp_io_sync_en_c2t  
	.stg2_db0_clk_stop_in_c2b ( stg2_db0_clk_stop_c1b  ),// UNDRIVEN stg2_db0_clk_stop_c2b  
	.stg2_dmu_io_clk_stop_in_c2b ( stg2_dmu_io_clk_stop_c1b  ), // UNDRIVEN stg2_dmu_io_clk_stop_c2b  
	.stg2_dmu_peu_por_in_c2b ( stg2_dmu_peu_por_c1b  ), // UNDRIVEN stg2_dmu_peu_por_c2b  
	.stg2_dmu_peu_wmr_in_c2b ( stg2_dmu_peu_wmr_c1b  ), // UNDRIVEN stg2_dmu_peu_wmr_c2b  
	.stg2_dr_sync_en_in_c2t ( stg2_dr_sync_en_c1t  ),// stg2_dr_sync_en_c2t  UNDRIVEN 
	.stg2_io_cmp_sync_en_in_c2b ( stg2_io_cmp_sync_en_c1b  ),// UNDRIVEN stg2_io_cmp_sync_en_c2b  
	.stg2_io_cmp_sync_en_in_c2t ( stg2_io_cmp_sync_en_c1t  ),// UNDRIVEN stg2_io_cmp_sync_en_c2t  
	.stg2_io_out_in_c2t ( stg2_io_out_c1t  ),// UNDRIVEN stg2_io_out_c2t  
	.stg2_io_out_in_c2b ( stg2_io_out_c1b  ),// UNDRIVEN stg2_io_out_c2b  
	.stg2_l2_por_in_c2b ( stg2_l2_por_c1b  ),// UNDRIVEN stg2_l2_por_c2b  
	.stg2_l2_por_in_c2t ( stg2_l2_por_c1t  ),// UNDRIVEN stg2_l2_por_c2t  
	.stg2_l2_wmr_in_c2b ( stg2_l2_wmr_c1b  ),// UNDRIVEN stg2_l2_wmr_c2b  
	.stg2_l2_wmr_in_c2t ( stg2_l2_wmr_c1t  ),// UNDRIVEN stg2_l2_wmr_c2t  
	.stg2_l2b0_clk_stop_in_c2t ( stg2_l2b0_clk_stop_c1t  ), // UNDRIVEN stg2_l2b0_clk_stop_c2t 
	.stg2_l2b1_clk_stop_in_c2t ( stg2_l2b1_clk_stop_c1t  ), // UNDRIVEN stg2_l2b1_clk_stop_c2t  
	.stg2_l2b2_clk_stop_in_c2b ( stg2_l2b2_clk_stop_c1b  ),// UNDRIVEN stg2_l2b2_clk_stop_c2b  
	.stg2_l2b3_clk_stop_in_c2b ( stg2_l2b3_clk_stop_c1b  ),// UNDRIVEN stg2_l2b3_clk_stop_c2b  
	.stg2_l2d0_clk_stop_in_c2t ( stg2_l2d0_clk_stop_c1t  ),// UNDRIVEN stg2_l2d0_clk_stop_c2t  
	.stg2_l2d1_clk_stop_in_c2t ( stg2_l2d1_clk_stop_c1t  ),// UNDRIVEN stg2_l2d1_clk_stop_c2t  
	.stg2_l2d2_clk_stop_in_c2b ( stg2_l2d2_clk_stop_c1b  ),// UNDRIVEN stg2_l2d2_clk_stop_c2b  
	.stg2_l2d3_clk_stop_in_c2b ( stg2_l2d3_clk_stop_c1b  ),// UNDRIVEN stg2_l2d3_clk_stop_c2b  
	.stg2_l2t0_clk_stop_in_c2t ( stg2_l2t0_clk_stop_c1t  ),// UNDRIVEN stg2_l2t0_clk_stop_c2t  
	.stg2_l2t1_clk_stop_in_c2t ( stg2_l2t1_clk_stop_c1t  ),// UNDRIVEN stg2_l2t1_clk_stop_c2t  
	.stg2_l2t2_clk_stop_in_c2b ( stg2_l2t2_clk_stop_c1b  ),// UNDRIVEN stg2_l2t2_clk_stop_c2b  
	.stg2_l2t3_clk_stop_in_c2bz ( stg2_l2t3_clk_stop_c1b  ),// UNDRIVEN stg2_l2t3_clk_stop_c2bz  
	.stg2_l2t5_clk_stop_in_c2t ( stg2_l2t5_clk_stop_c1t  ),// UNDRIVEN stg2_l2t5_clk_stop_c2t  
	.stg2_l2t7_clk_stop_in_c2b ( stg2_l2t7_clk_stop_c1b  ),// UNDRIVEN stg2_l2t7_clk_stop_c2b  
	.stg2_mio_io2x_sync_en_in_c2t ( stg2_mio_io2x_sync_en_c1t  ), // UNDRIVEN stg2_mio_io2x_sync_en_c2t  
	.stg2_mio_clk_stop_in_c2t ( stg2_mio_clk_stop_c1t ),// UNDRIVEN stg2_mio_clk_stop_c2t 
	.stg2_ncu_clk_stop_in_c2b ( stg2_ncu_clk_stop_c1b  ),// UNDRIVEN stg2_ncu_clk_stop_c2b  
	.stg2_ncu_io_clk_stop_in_c2b ( stg2_ncu_io_clk_stop_c1b  ), // UNDRIVEN stg2_ncu_io_clk_stop_c2b  
	.stg2_peu_io_clk_stop_in_c2b ( stg2_peu_io_clk_stop_c1b  ), // UNDRIVEN stg2_peu_io_clk_stop_c2b  
	.stg2_sii_clk_stop_in_c2b ( stg2_sii_clk_stop_c1b  ), // UNDRIVEN stg2_sii_clk_stop_c2b  
	.stg2_sii_io_clk_stop_in_c2b ( stg2_sii_io_clk_stop_c1b  ), // UNDRIVEN stg2_sii_io_clk_stop_c2b  
	.stg2_spc0_clk_stop_in_c2t ( stg2_spc0_clk_stop_c1t  ), // UNDRIVEN stg2_spc0_clk_stop_c2t  
	.stg2_spc1_clk_stop_in_c2t ( stg2_spc1_clk_stop_c1t  ), // UNDRIVEN stg2_spc1_clk_stop_c2t  
	.stg2_spc2_clk_stop_in_c2b ( stg2_spc2_clk_stop_c1b  ), // UNDRIVEN stg2_spc2_clk_stop_c2b  
	.stg2_spc3_clk_stop_in_c2b ( stg2_spc3_clk_stop_c1b  ), // UNDRIVEN stg2_spc3_clk_stop_c2b  
	.stg2_spc5_clk_stop_in_c2t ( stg2_spc5_clk_stop_c1t  ), // UNDRIVEN stg2_spc5_clk_stop_c2t  
	.stg2_spc7_clk_stop_in_c2b ( stg2_spc7_clk_stop_c1b  ), // UNDRIVEN stg2_spc7_clk_stop_c2b  
    .stg2_io2x_sync_en_in_c2t  ( 1'b0 ), // ERROR: stg2_mio_io2x_sync_en_c2t 
	.stg3_ccx_clk_stop_in_c2b ( stg3_ccx_clk_stop_c2b  ),
	.stg3_cmp_io_sync_en_in_c2b ( stg3_cmp_io_sync_en_c2b  ), // CHECK
	.stg3_cmp_io_sync_en_in_c2t ( stg3_cmp_io_sync_en_c2t  ), // CHECK
	.stg3_cmp_io_sync_en_in_c3b ( stg3_cmp_io_sync_en_c2b  ),// UNDRIVEN stg3_cmp_io_sync_en_c3b  
	.stg3_cmp_io_sync_en_in_c3t ( stg3_cmp_io_sync_en_c2t  ),// UNDRIVEN stg3_cmp_io_sync_en_c3t  
	.stg3_db0_clk_stop_in_c3b ( stg3_db0_clk_stop_c2b  ),// UNDRIVEN stg3_db0_clk_stop_c3b  
	.stg3_dmu_io_clk_stop_in_c3b ( stg3_dmu_io_clk_stop_c2b  ),// UNDRIVEN stg3_dmu_io_clk_stop_c3b  
	.stg3_dmu_peu_por_in_c3b ( stg3_dmu_peu_por_c2b  ), // UNDRIVEN stg3_dmu_peu_por_c3b  
	.stg3_dmu_peu_wmr_in_c3b ( stg3_dmu_peu_wmr_c2b  ), // UNDRIVEN stg3_dmu_peu_wmr_c3b  
	.stg3_dr_sync_en_in_c3t ( stg3_dr_sync_en_c2t  ),	// stg3_dr_sync_en_c3t   UNDRIVEN
	.stg3_io2x_sync_en_in_c2t ( stg3_mio_io2x_sync_en_c2t ), // UNDRIVEN stg3_io2x_sync_en_c2t  
	.stg3_io_cmp_sync_en_in_c2b ( stg3_io_cmp_sync_en_c2b  ), // CHECK
	.stg3_io_cmp_sync_en_in_c2t ( stg3_io_cmp_sync_en_c2t  ), // CHECK
	.stg3_io_cmp_sync_en_in_c3b ( stg3_io_cmp_sync_en_c2b  ), // UNDRIVEN stg3_io_cmp_sync_en_c3b  
	.stg3_io_cmp_sync_en_in_c3t ( stg3_io_cmp_sync_en_c2t  ), // UNDRIVEN stg3_io_cmp_sync_en_c3t  
	.stg3_io_out_in_c3b ( stg3_io_out_c2b  ), // UNDRIVEN stg3_io_out_c3b  
	.stg3_io_out_in_c3t ( stg3_io_out_c2t  ), // UNDRIVEN stg3_io_out_c3t  
	.stg3_l2_por_in_c2b ( stg3_l2_por_c2b  ),
	.stg3_l2_por_in_c2t ( stg3_l2_por_c2t  ),
	.stg3_l2_por_in_c3b ( stg3_l2_por_c2b  ), // UNDRIVEN stg3_l2_por_c3b  
	.stg3_l2_por_in_c3t ( stg3_l2_por_c2t  ), // UNDRIVEN stg3_l2_por_c3t  
	.stg3_l2_wmr_in_c2b ( stg3_l2_wmr_c2b  ),
	.stg3_l2_wmr_in_c2t ( stg3_l2_wmr_c2t  ),
	.stg3_l2_wmr_in_c3b ( stg3_l2_wmr_c2b  ), // UNDRIVEN stg3_l2_wmr_c3b  
	.stg3_l2_wmr_in_c3t ( stg3_l2_wmr_c2t  ), // UNDRIVEN stg3_l2_wmr_c3t  
	.stg3_l2b0_clk_stop_in_c3t ( stg3_l2b0_clk_stop_c2t  ), // UNDRIVEN stg3_l2b0_clk_stop_c3t  
	.stg3_l2b1_clk_stop_in_c3t ( stg3_l2b1_clk_stop_c2t  ), // UNDRIVEN stg3_l2b1_clk_stop_c3t  
	.stg3_l2b2_clk_stop_in_c3b ( stg3_l2b2_clk_stop_c2b  ), // UNDRIVEN stg3_l2b2_clk_stop_c3b  
	.stg3_l2b3_clk_stop_in_c3b ( stg3_l2b3_clk_stop_c2b  ), // UNDRIVEN stg3_l2b3_clk_stop_c3b  
	.stg3_l2d0_clk_stop_in_c3t ( stg3_l2d0_clk_stop_c2t  ), // UNDRIVEN stg3_l2d0_clk_stop_c3t  
	.stg3_l2d1_clk_stop_in_c3t ( stg3_l2d1_clk_stop_c2t  ), // UNDRIVEN stg3_l2d1_clk_stop_c3t  
	.stg3_l2d2_clk_stop_in_c3b ( stg3_l2d2_clk_stop_c2b  ), // UNDRIVEN stg3_l2d2_clk_stop_c3b  
	.stg3_l2d3_clk_stop_in_c3b ( stg3_l2d3_clk_stop_c2b  ), // UNDRIVEN stg3_l2d3_clk_stop_c3b  
	.stg3_l2t0_clk_stop_in_c3t ( stg3_l2t0_clk_stop_c2t  ), // UNDRIVEN stg3_l2t0_clk_stop_c3t  
	.stg3_l2t1_clk_stop_in_c2t ( stg3_l2t1_clk_stop_c2t  ), // UNDRIVEN stg3_l2t1_clk_stop_c2t  
	.stg3_l2t2_clk_stop_in_c3b ( stg3_l2t2_clk_stop_c2b  ), // UNDRIVEN stg3_l2t2_clk_stop_c3b  
	.stg3_l2t3_clk_stop_in_c2b ( stg3_l2t3_clk_stop_c2b  ),
	.stg3_l2t5_clk_stop_in_c2t ( stg3_l2t5_clk_stop_c2t  ),
	.stg3_l2t7_clk_stop_in_c2b ( stg3_l2t7_clk_stop_c2b  ),
	.stg3_mcu0_clk_stop_in_c3t ( stg3_mcu0_clk_stop_c2t  ), // UNDRIVEN stg3_mcu0_clk_stop_c3t  
	.stg2_mcu0_dr_clk_stop_in_c4t ( stg2_mcu0_dr_clk_stop_c2b  ), // UNDRIVEN stg2_mcu0_dr_clk_stop_c3t  
	.stg3_mcu0_io_clk_stop_in_c3t ( stg3_mcu0_io_clk_stop_c2t  ), // UNDRIVEN stg3_mcu0_io_clk_stop_c3t  
	.stg3_mcu1_clk_stop_in_c3t ( stg3_mcu1_clk_stop_c2t  ), // UNDRIVEN stg3_mcu1_clk_stop_c3t  
	.stg2_mcu1_dr_clk_stop_in_c4t ( stg2_mcu1_dr_clk_stop_c2b ), // UD stg2_mcu1_dr_clk_stop_c3t  
	.stg3_mcu1_io_clk_stop_in_c3t ( stg3_mcu1_io_clk_stop_c2t ), // UD stg3_mcu1_io_clk_stop_c3t  
	.stg3_mio_clk_stop_in_c2t ( stg3_mio_clk_stop_c2t  ),
	.stg3_mio_clk_stop_in_c3t ( stg3_mio_clk_stop_c2t  ), // UNDRIVEN stg3_mio_clk_stop_c3t  
	.stg3_mio_io2x_sync_en_in_c3t ( stg3_mio_io2x_sync_en_c2t  ),// UNDRIVEN stg3_mio_io2x_sync_en_c3t  
	.stg3_ncu_clk_stop_in_c3b ( stg3_ncu_clk_stop_c2b  ),	// UNDRIVEN stg3_ncu_clk_stop_c3b  
	.stg3_ncu_io_clk_stop_in_c3b ( stg3_ncu_io_clk_stop_c2b  ),// UNDRIVEN stg3_ncu_io_clk_stop_c3b  
	.stg3_peu_io_clk_stop_in_c3b ( stg3_peu_io_clk_stop_c2b  ),// UNDRIVEN stg3_peu_io_clk_stop_c3b  
	.stg3_sii_clk_stop_in_c3b ( stg3_sii_clk_stop_c2b  ),// UNDRIVEN stg3_sii_clk_stop_c3b  
	.stg3_sii_io_clk_stop_in_c3b ( stg3_sii_io_clk_stop_c2b  ),// UNDRIVEN stg3_sii_io_clk_stop_c3b  
	.stg3_spc0_clk_stop_in_c3t ( stg3_spc0_clk_stop_c2t  ),	// UNDRIVEN stg3_spc0_clk_stop_c3t  
	.stg3_spc1_clk_stop_in_c2t ( stg3_spc1_clk_stop_c2t  ),	// UNDRIVEN stg3_spc1_clk_stop_c2b  
	.stg3_spc2_clk_stop_in_c3b ( stg3_spc2_clk_stop_c2b  ), // UNDRIVEN stg3_spc2_clk_stop_c3b  
	.stg3_spc3_clk_stop_in_c2b ( stg3_spc3_clk_stop_c2b ),		
	.stg3_spc5_clk_stop_in_c2t ( stg3_spc5_clk_stop_c2t  ), // UNDRIVEN stg3_spc5_clk_stop_c2b  
	.stg3_spc7_clk_stop_in_c2b ( stg3_spc7_clk_stop_c2b ),		
	.stg4_cmp_io_sync_en_in_c3b ( stg4_cmp_io_sync_en_c3b  ),
	.stg4_cmp_io_sync_en_in_c3t ( stg4_cmp_io_sync_en_c3t  ),
	.stg4_db0_clk_stop_c3b ( stg4_db0_clk_stop_c3b ),		// ERROR!! should be stg4_db0_clk_stop_in_c3b 
	.stg4_dmu_io_clk_stop_in_c3b ( stg4_dmu_io_clk_stop_c3b  ),
	.stg4_dmu_peu_por_in_c3b ( stg4_dmu_peu_por_c3b  ),
	.stg4_dmu_peu_wmr_in_c3b ( stg4_dmu_peu_wmr_c3b  ),
	.stg4_dr_sync_en_in_c3t ( stg4_dr_sync_en_c3t  ),
	.stg4_io2x_sync_en_in_c3t ( stg4_mio_io2x_sync_en_c3t ), // UNDRIVEN stg4_io2x_sync_en_c3t 
	.stg4_io_cmp_sync_en_in_c3b ( stg4_io_cmp_sync_en_c3b  ),
	.stg4_io_cmp_sync_en_in_c3t ( stg4_io_cmp_sync_en_c3t  ),
	.stg4_io_out_in_c3b ( stg4_io_out_c3b  ),
	.stg4_io_out_in_c3t ( stg4_io_out_c3t  ),
	.stg4_l2_por_in_c3b ( stg4_l2_por_c3b  ),
	.stg4_l2_por_in_c3t ( stg4_l2_por_c3t  ),
	.stg4_l2_wmr_in_c3b ( stg4_l2_wmr_c3b  ),
	.stg4_l2_wmr_in_c3t ( stg4_l2_wmr_c3t  ),
	.stg4_l2b0_clk_stop_in_c3t ( stg4_l2b0_clk_stop_c3t  ),
	.stg4_l2b1_clk_stop_in_c3t ( stg4_l2b1_clk_stop_c3t  ),
	.stg4_l2b2_clk_stop_in_c3b ( stg4_l2b2_clk_stop_c3b  ),
	.stg4_l2b3_clk_stop_in_c3b ( stg4_l2b3_clk_stop_c3b  ),
	.stg4_l2d0_clk_stop_in_c3t ( stg4_l2d0_clk_stop_c3t  ),
	.stg4_l2d1_clk_stop_in_c3t ( stg4_l2d1_clk_stop_c3t  ),
	.stg4_l2d2_clk_stop_in_c3b ( stg4_l2d2_clk_stop_c3b  ),
	.stg4_l2d3_clk_stop_in_c3b ( stg4_l2d3_clk_stop_c3b  ),
	.stg4_l2t0_clk_stop_in_c3t ( stg4_l2t0_clk_stop_c3t  ),
	.stg4_l2t2_clk_stop_in_c3b ( stg4_l2t2_clk_stop_c3b  ),
//	.stg4_mcu1_dr_clk_stop_in_c3t ( stg4_mcu1_dr_clk_stop_c3t  ),
	.stg4_mcu0_clk_stop_in_c3t ( stg4_mcu0_clk_stop_c3t  ),
//	.stg4_mcu0_dr_clk_stop_in_c3t ( stg4_mcu0_dr_clk_stop_c3t  ),
	.stg4_mcu0_io_clk_stop_in_c3t ( stg4_mcu0_io_clk_stop_c3t  ),
	.stg4_mcu1_clk_stop_in_c3t ( stg4_mcu1_clk_stop_c3t  ),
	.stg4_mcu1_io_clk_stop_in_c3t ( stg4_mcu1_io_clk_stop_c3t  ),
	.stg4_mio_clk_stop_in_c3t ( stg4_mio_clk_stop_c3t  ), // UNDRIVEN stg4_mio_clk_stop_c3tz  
	.stg4_ncu_clk_stop_in_c3b ( stg4_ncu_clk_stop_c3b  ),
	.stg4_ncu_io_clk_stop_c3b ( stg4_ncu_io_clk_stop_c3b ),		// ERROR!! - should be stg4_ncu_io_clk_stop_in_c3b 
	.stg4_peu_io_clk_stop_in_c3b ( stg4_peu_io_clk_stop_c3b  ),
	.stg4_sii_clk_stop_in_c3b ( stg4_sii_clk_stop_c3b  ),
	.stg4_sii_io_clk_stop_in_c3b ( stg4_sii_io_clk_stop_c3b  ),
	.stg4_spc0_clk_stop_in_c3t ( stg4_spc0_clk_stop_c3t  ),
	.stg4_spc2_clk_stop_in_c3b ( stg4_spc2_clk_stop_c3b  ),
	.stg2_mcu0_io_clk_stop_in_c2t ( stg2_mcu0_io_clk_stop_c1t ), // UD stg2_mcu0_io_clk_stop_c2t 
//	.stg2_mcu0_dr_clk_stop_in_c2t ( stg2_mcu0_dr_clk_stop_c1t ), // UD stg2_mcu0_dr_clk_stop_c2t 
//	.stg2_mcu1_dr_clk_stop_in_c2t ( stg2_mcu1_dr_clk_stop_c1t ), // UD stg2_mcu1_dr_clk_stop_c2t 
	.stg2_mcu1_io_clk_stop_in_c2t ( stg2_mcu1_io_clk_stop_c1t ), // UD stg2_mcu1_io_clk_stop_c2t 

	// STAGED OUTPUTS
//	.stg3_mcu0_dr_clk_stop_out_c2t ( stg3_mcu0_dr_clk_stop_c2t ),
	.stg3_mcu0_io_clk_stop_out_c2t ( stg3_mcu0_io_clk_stop_c2t ),
//	.stg3_mcu1_dr_clk_stop_out_c2t ( stg3_mcu1_dr_clk_stop_c2t ),
	.stg3_mcu1_io_clk_stop_out_c2t ( stg3_mcu1_io_clk_stop_c2t ),
	.stg1_ccx_clk_stop_out_c1b ( stg1_ccx_clk_stop_c1b  ),
	.stg1_cmp_io_sync_en_out_c1b ( stg1_cmp_io_sync_en_c1b  ),
	.stg1_cmp_io_sync_en_out_c1t ( stg1_cmp_io_sync_en_c1t  ),
	.stg1_db0_clk_stop_out_c1b ( stg1_db0_clk_stop_c1b  ),
	.stg1_dmu_io_clk_stop_out_c1b ( stg1_dmu_io_clk_stop_c1b  ),
	.stg1_dmu_peu_por_out_c1b ( stg1_dmu_peu_por_c1b  ),
	.stg1_dmu_peu_wmr_out_c1b ( stg1_dmu_peu_wmr_c1b  ),
	.stg1_dr_sync_en_out_c1t ( stg1_dr_sync_en_c1t  ),
	.stg1_io2x_out_out_c1b ( stg1_io2x_out_c1b  ),
	.stg1_io2x_sync_en_out_c1b ( stg1_io2x_sync_en_c1b  ),
	.stg1_io2x_sync_en_out_c1t ( stg1_io2x_sync_en_c1t  ),
	.stg1_io_cmp_sync_en_out_c1b ( stg1_io_cmp_sync_en_c1b  ),
	.stg1_io_cmp_sync_en_out_c1t ( stg1_io_cmp_sync_en_c1t  ),
	.stg1_io_out_out_c1b ( stg1_io_out_c1b  ),
	.stg1_io_out_out_c1t ( stg1_io_out_c1t  ),
	.stg1_l2b0_clk_stop_out_c1t ( stg1_l2b0_clk_stop_c1t  ),
	.stg1_l2b1_clk_stop_out_c1t ( stg1_l2b1_clk_stop_c1t  ),
	.stg1_l2b2_clk_stop_out_c1b ( stg1_l2b2_clk_stop_c1b  ),
	.stg1_l2b3_clk_stop_out_c1b ( stg1_l2b3_clk_stop_c1b  ),
	.stg1_l2b4_clk_stop_out_c1t ( stg1_l2b4_clk_stop_c1t  ),
	.stg1_l2b5_clk_stop_out_c1t ( stg1_l2b5_clk_stop_c1t  ),
	.stg1_l2d0_clk_stop_out_c1t ( stg1_l2d0_clk_stop_c1t  ),
	.stg1_l2d1_clk_stop_out_c1t ( stg1_l2d1_clk_stop_c1t  ),
	.stg1_l2d2_clk_stop_out_c1b ( stg1_l2d2_clk_stop_c1b  ),
	.stg1_l2d3_clk_stop_out_c1b ( stg1_l2d3_clk_stop_c1b  ),
	.stg1_l2d4_clk_stop_out_c1t ( stg1_l2d4_clk_stop_c1t  ),
	.stg1_l2d5_clk_stop_out_c1t ( stg1_l2d5_clk_stop_c1t  ),
//	.stg1_l2d6_clk_stop_out_c1b ( stg1_l2d6_clk_stop_c1b  ),  // ECO1.1 -mh157021
	.stg1_l2d7_clk_stop_out_c1b ( stg1_l2d7_clk_stop_c1b  ),  // ECO1.1 -mh157021
	.stg1_l2t0_clk_stop_out_c1t ( stg1_l2t0_clk_stop_c1t  ),
	.stg1_l2t1_clk_stop_out_c1t ( stg1_l2t1_clk_stop_c1t  ),
	.stg1_l2t2_clk_stop_out_c1b ( stg1_l2t2_clk_stop_c1b  ),
	.stg1_l2t3_clk_stop_out_c1b ( stg1_l2t3_clk_stop_c1b  ),
	.stg1_l2t5_clk_stop_out_c1t ( stg1_l2t5_clk_stop_c1t  ),
	.stg1_l2t7_clk_stop_out_c1b ( stg1_l2t7_clk_stop_c1b  ),
	.stg1_mac_io_clk_stop_out_c1b ( stg1_mac_io_clk_stop_c1b  ),
	.stg1_mcu0_clk_stop_out_c1t ( stg1_mcu0_clk_stop_c1t  ),
	.stg1_mcu0_dr_clk_stop_out_c1t ( stg1_mcu0_dr_clk_stop_c1t  ),
	.stg1_mcu0_io_clk_stop_out_c1t ( stg1_mcu0_io_clk_stop_c1t  ),
	.stg1_mcu1_clk_stop_out_c1t ( stg1_mcu1_clk_stop_c1t  ),
	.stg1_mcu1_dr_clk_stop_out_c1t ( stg1_mcu1_dr_clk_stop_c1t  ),
	.stg1_mcu1_io_clk_stop_out_c1t ( stg1_mcu1_io_clk_stop_c1t  ),
	.stg1_mio_clk_stop_out_c1t ( stg1_mio_clk_stop_c1t  ),
	.stg3_mio_clk_stop_out_c2t ( stg3_mio_clk_stop_c2t  ),
	.stg1_ncu_clk_stop_out_c1b ( stg1_ncu_clk_stop_c1b  ),
	.stg1_ncu_io_clk_stop_out_c1b ( stg1_ncu_io_clk_stop_c1b  ),
	.stg1_peu_io_clk_stop_out_c1b ( stg1_peu_io_clk_stop_c1b  ),
	.stg1_rdp_io_clk_stop_out_c1b ( stg1_rdp_io_clk_stop_c1b  ),
	.stg1_rst_l2_por_out_c1b ( stg1_rst_l2_por_c1b  ),
	.stg1_rst_l2_por_out_c1t ( stg1_rst_l2_por_c1t  ),
	.stg1_rst_l2_wmr_out_c1b ( stg1_rst_l2_wmr_c1b  ),
	.stg1_rst_l2_wmr_out_c1t ( stg1_rst_l2_wmr_c1t  ),
	.stg1_rst_niu_mac_out_c1b ( stg1_rst_niu_mac_c1b  ),
	.stg1_rst_niu_wmr_out_c1b ( stg1_rst_niu_wmr_c1b  ),
	.stg1_rtx_io_clk_stop_out_c1b ( stg1_rtx_io_clk_stop_c1b  ),
	.stg1_sii_clk_stop_out_c1b ( stg1_sii_clk_stop_c1b  ),
	.stg1_sii_io_clk_stop_out_c1b ( stg1_sii_io_clk_stop_c1b  ),
	.stg1_spc0_clk_stop_out_c1t ( stg1_spc0_clk_stop_c1t  ),
	.stg1_spc1_clk_stop_out_c1t ( stg1_spc1_clk_stop_c1t  ),
	.stg1_spc2_clk_stop_out_c1b ( stg1_spc2_clk_stop_c1b  ),
	.stg1_spc3_clk_stop_out_c1b ( stg1_spc3_clk_stop_c1b  ),
	.stg1_spc4_clk_stop_out_c1t ( stg1_spc4_clk_stop_c1t  ),
	.stg1_spc5_clk_stop_out_c1t ( stg1_spc5_clk_stop_c1t  ),
	.stg1_spc6_clk_stop_out_c1b ( stg1_spc6_clk_stop_c1b  ),
	.stg1_spc7_clk_stop_out_c1b ( stg1_spc7_clk_stop_c1b  ),
	.stg1_tds_io_clk_stop_out_c1b ( stg1_tds_io_clk_stop_c1b  ),
	.stg2_ccx_clk_stop_out_c1b ( stg2_ccx_clk_stop_c1b  ),
	.stg2_cmp_io_sync_en_out_c1b ( stg2_cmp_io_sync_en_c1b  ),
	.stg2_cmp_io_sync_en_out_c1t ( stg2_cmp_io_sync_en_c1t  ),
	.stg2_db0_clk_stop_out_c1b ( stg2_db0_clk_stop_c1b  ),
	.stg2_dmu_io_clk_stop_out_c1b ( stg2_dmu_io_clk_stop_c1b  ),
	.stg2_dmu_peu_por_out_c1b ( stg2_dmu_peu_por_c1b  ),
	.stg2_dmu_peu_wmr_out_c1b ( stg2_dmu_peu_wmr_c1b  ),
	.stg2_dr_sync_en_out_c1t ( stg2_dr_sync_en_c1t  ),
	.stg2_io_cmp_sync_en_out_c1b ( stg2_io_cmp_sync_en_c1b  ),
	.stg2_io_cmp_sync_en_out_c1t ( stg2_io_cmp_sync_en_c1t  ),
	.stg2_io_out_out_c1t ( stg2_io_out_c1t  ),
	.stg2_io_out_out_c1b ( stg2_io_out_c1b  ), // marked
	.stg2_l2_por_out_c1b ( stg2_l2_por_c1b  ),
	.stg2_l2_por_out_c1t ( stg2_l2_por_c1t  ),
	.stg2_l2_wmr_out_c1b ( stg2_l2_wmr_c1b  ),
	.stg2_l2_wmr_out_c1t ( stg2_l2_wmr_c1t  ),
	.stg2_l2b0_clk_stop_out_c1t ( stg2_l2b0_clk_stop_c1t  ),
	.stg2_l2b1_clk_stop_out_c1t ( stg2_l2b1_clk_stop_c1t  ),
	.stg2_l2b2_clk_stop_out_c1b ( stg2_l2b2_clk_stop_c1b  ),
	.stg2_l2b3_clk_stop_out_c1b ( stg2_l2b3_clk_stop_c1b  ),
	.stg2_l2d0_clk_stop_out_c1t ( stg2_l2d0_clk_stop_c1t  ),
	.stg2_l2d1_clk_stop_out_c1t ( stg2_l2d1_clk_stop_c1t  ),
	.stg2_l2d2_clk_stop_out_c1b ( stg2_l2d2_clk_stop_c1b  ),
	.stg2_l2d3_clk_stop_out_c1b ( stg2_l2d3_clk_stop_c1b  ),
	.stg2_l2t0_clk_stop_out_c1t ( stg2_l2t0_clk_stop_c1t  ),
	.stg2_l2t1_clk_stop_out_c1t ( stg2_l2t1_clk_stop_c1t  ),
	.stg2_l2t2_clk_stop_out_c1b ( stg2_l2t2_clk_stop_c1b  ),
	.stg2_l2t3_clk_stop_out_c1b ( stg2_l2t3_clk_stop_c1b  ),
	.stg2_l2t5_clk_stop_out_c1t ( stg2_l2t5_clk_stop_c1t  ),
	.stg2_l2t7_clk_stop_out_c1b ( stg2_l2t7_clk_stop_c1b  ),
	.stg2_mcu0_clk_stop_out_c1t ( stg2_mcu0_clk_stop_c1t  ),
	.stg2_mcu0_dr_clk_stop_out_c2b ( stg2_mcu0_dr_clk_stop_c2b  ),
	.stg2_mcu1_dr_clk_stop_out_c2b ( stg2_mcu1_dr_clk_stop_c2b  ),
	.stg2_mcu0_io_clk_stop_out_c1t ( stg2_mcu0_io_clk_stop_c1t  ),
	.stg2_mcu1_clk_stop_out_c1t ( stg2_mcu1_clk_stop_c1t  ),
	.stg2_mcu1_io_clk_stop_out_c1t ( stg2_mcu1_io_clk_stop_c1t  ),
	.stg2_mio_clk_stop_out_c1t ( stg2_mio_clk_stop_c1t  ),
	.stg2_mio_io2x_sync_en_out_c1t ( stg2_mio_io2x_sync_en_c1t  ),
//     .stg2_mio_io2x_sync_en_out_c2t  (stg2_mio_io2x_sync_en_c2t ),
	.stg2_ncu_clk_stop_out_c1b ( stg2_ncu_clk_stop_c1b  ),
	.stg2_ncu_io_clk_stop_out_c1b ( stg2_ncu_io_clk_stop_c1b  ),
	.stg2_peu_io_clk_stop_out_c1b ( stg2_peu_io_clk_stop_c1b  ),
	.stg2_sii_clk_stop_out_c1b ( stg2_sii_clk_stop_c1b  ),
	.stg2_sii_io_clk_stop_out_c1b ( stg2_sii_io_clk_stop_c1b  ),
	.stg2_spc0_clk_stop_out_c1t ( stg2_spc0_clk_stop_c1t  ),
	.stg2_spc1_clk_stop_out_c1t ( stg2_spc1_clk_stop_c1t  ),
	.stg2_spc2_clk_stop_out_c1b ( stg2_spc2_clk_stop_c1b  ),
	.stg2_spc3_clk_stop_out_c1b ( stg2_spc3_clk_stop_c1b  ),
	.stg2_spc5_clk_stop_out_c1t ( stg2_spc5_clk_stop_c1t  ),
	.stg2_spc7_clk_stop_out_c1b ( stg2_spc7_clk_stop_c1b  ),
	.stg3_ccx_clk_stop_out_c2b ( stg3_ccx_clk_stop_c2b  ),
	.stg3_cmp_io_sync_en_out_c2b ( stg3_cmp_io_sync_en_c2b  ),
	.stg3_cmp_io_sync_en_out_c2t ( stg3_cmp_io_sync_en_c2t  ),
	.stg3_db0_clk_stop_out_c2b ( stg3_db0_clk_stop_c2b  ),
	.stg3_dmu_io_clk_stop_out_c2b ( stg3_dmu_io_clk_stop_c2b  ),
	.stg3_dmu_peu_por_out_c2b ( stg3_dmu_peu_por_c2b  ),
	.stg3_dmu_peu_wmr_out_c2b ( stg3_dmu_peu_wmr_c2b  ),
	.stg3_dr_sync_en_out_c2t ( stg3_dr_sync_en_c2t  ),
	.stg3_io_cmp_sync_en_out_c2b ( stg3_io_cmp_sync_en_c2b  ),
	.stg3_io_cmp_sync_en_out_c2t ( stg3_io_cmp_sync_en_c2t  ),
	.stg3_io_out_out_c2t ( stg3_io_out_c2t  ),
	.stg3_l2_por_out_c2b ( stg3_l2_por_c2b  ),
	.stg3_l2_por_out_c2t ( stg3_l2_por_c2t  ),
	.stg3_l2_wmr_out_c2b ( stg3_l2_wmr_c2b  ),
	.stg3_l2_wmr_out_c2t ( stg3_l2_wmr_c2t  ),
	.stg3_l2b0_clk_stop_out_c2t ( stg3_l2b0_clk_stop_c2t  ),
	.stg3_l2b1_clk_stop_out_c2t ( stg3_l2b1_clk_stop_c2t  ),
	.stg3_l2b2_clk_stop_out_c2b ( stg3_l2b2_clk_stop_c2b  ),
	.stg3_l2b3_clk_stop_out_c2b ( stg3_l2b3_clk_stop_c2b  ),
	.stg3_l2d0_clk_stop_out_c2t ( stg3_l2d0_clk_stop_c2t  ),
	.stg3_l2d1_clk_stop_out_c2t ( stg3_l2d1_clk_stop_c2t  ),
	.stg3_l2d2_clk_stop_out_c2b ( stg3_l2d2_clk_stop_c2b  ),
	.stg3_l2d3_clk_stop_out_c2b ( stg3_l2d3_clk_stop_c2b  ),
	.stg3_l2t0_clk_stop_out_c2t ( stg3_l2t0_clk_stop_c2t  ),
	.stg3_l2t1_clk_stop_out_c2t ( stg3_l2t1_clk_stop_c2t  ),
	.stg3_l2t2_clk_stop_out_c2b ( stg3_l2t2_clk_stop_c2b  ),
	.stg3_l2t3_clk_stop_out_c2b ( stg3_l2t3_clk_stop_c2b  ),
	.stg3_l2t5_clk_stop_out_c2t ( stg3_l2t5_clk_stop_c2t  ),
	.stg3_l2t7_clk_stop_out_c2b ( stg3_l2t7_clk_stop_c2b  ),
	.stg3_mio_io2x_sync_en_out_c2t ( stg3_mio_io2x_sync_en_c2t  ),
//	.stg3_mcu0_dr_clk_stop_out_c2t ( stg3_mcu0_dr_clk_stop_c2t  ),
//	.stg3_mcu1_dr_clk_stop_out_c2t ( stg3_mcu1_dr_clk_stop_c2t  ),
	.stg3_ncu_clk_stop_out_c2b ( stg3_ncu_clk_stop_c2b  ),
	.stg3_ncu_io_clk_stop_out_c2b ( stg3_ncu_io_clk_stop_c2b  ),
	.stg3_io_out_out_c2b ( stg3_io_out_c2b  ),	 // marked
	.stg3_peu_io_clk_stop_out_c2b ( stg3_peu_io_clk_stop_c2b  ),
	.stg3_sii_clk_stop_out_c2b ( stg3_sii_clk_stop_c2b  ),
	.stg3_sii_io_clk_stop_out_c2b ( stg3_sii_io_clk_stop_c2b  ),
	.stg3_spc0_clk_stop_out_c2t ( stg3_spc0_clk_stop_c2t  ),
	.stg3_spc1_clk_stop_out_c2t ( stg3_spc1_clk_stop_c2t  ),
	.stg3_spc2_clk_stop_out_c2b ( stg3_spc2_clk_stop_c2b  ),
	.stg3_spc3_clk_stop_out_c2b ( stg3_spc3_clk_stop_c2b  ),
	.stg3_spc5_clk_stop_out_c2t ( stg3_spc5_clk_stop_c2t  ),
	.stg3_spc7_clk_stop_out_c2b ( stg3_spc7_clk_stop_c2b  ),
	.stg4_io2x_sync_en_c3t ( stg4_mio_io2x_sync_en_c3t ),	 // ECO1.3 .( stg4_io2x_sync_en_c3t ) -mh157021
	.stg4_cmp_io_sync_en_out_c3b ( stg4_cmp_io_sync_en_c3b  ),
	.stg4_cmp_io_sync_en_out_c3t ( stg4_cmp_io_sync_en_c3t  ),
	.stg4_db0_clk_stop_out_c3b ( stg4_db0_clk_stop_c3b  ),
	.stg4_dmu_io_clk_stop_out_c3b ( stg4_dmu_io_clk_stop_c3b  ),
	.stg4_dmu_peu_por_out_c3b ( stg4_dmu_peu_por_c3b  ),
	.stg4_dmu_peu_wmr_out_c3b ( stg4_dmu_peu_wmr_c3b  ),
	.stg4_dr_sync_en_out_c3t ( stg4_dr_sync_en_c3t  ),
    .stg3_io2x_sync_en_out_c2t  (stg3_io2x_sync_en_c2t), // ERROR : UNUSED
	// .stg4_io2x_sync_en_out_c2b ( stg4_io2x_sync_en_c2b  ),
	.stg4_io_cmp_sync_en_out_c3b ( stg4_io_cmp_sync_en_c3b  ),
	.stg4_io_cmp_sync_en_out_c3t ( stg4_io_cmp_sync_en_c3t  ),
	.stg4_io_out_out_c3b ( stg4_io_out_c3b  ),
	.stg4_io_out_out_c3t ( stg4_io_out_c3t  ),
	.stg4_l2_por_out_c3b ( stg4_l2_por_c3b  ),
	.stg4_l2_por_out_c3t ( stg4_l2_por_c3t  ),
	.stg4_l2_wmr_out_c3b ( stg4_l2_wmr_c3b  ),
	.stg4_l2_wmr_out_c3t ( stg4_l2_wmr_c3t  ),
	.stg4_l2b0_clk_stop_out_c3t ( stg4_l2b0_clk_stop_c3t  ),
	.stg4_l2b1_clk_stop_out_c3t ( stg4_l2b1_clk_stop_c3t  ),
	.stg4_l2b2_clk_stop_out_c3b ( stg4_l2b2_clk_stop_c3b  ),
	.stg4_l2b3_clk_stop_out_c3b ( stg4_l2b3_clk_stop_c3b  ),
	.stg4_l2d0_clk_stop_out_c3t ( stg4_l2d0_clk_stop_c3t  ),
	.stg4_l2d1_clk_stop_out_c3t ( stg4_l2d1_clk_stop_c3t  ),
	.stg4_l2d2_clk_stop_out_c3b ( stg4_l2d2_clk_stop_c3b  ),
	.stg4_l2d3_clk_stop_out_c3b ( stg4_l2d3_clk_stop_c3b  ),
	.stg4_l2t0_clk_stop_out_c3t ( stg4_l2t0_clk_stop_c3t  ),
	.stg4_l2t2_clk_stop_out_c3b ( stg4_l2t2_clk_stop_c3b  ),
	.stg4_mcu0_clk_stop_out_c3t ( stg4_mcu0_clk_stop_c3t  ),
//	.stg4_mcu0_dr_clk_stop_out_c3t ( stg4_mcu0_dr_clk_stop_c3t  ),
	.stg4_mcu0_io_clk_stop_out_c3t ( stg4_mcu0_io_clk_stop_c3t  ),
	.stg4_mcu1_clk_stop_out_c3t ( stg4_mcu1_clk_stop_c3t  ),
//	.stg4_mcu1_dr_clk_stop_out_c3t ( stg4_mcu1_dr_clk_stop_c3t  ),
	.stg4_mcu1_io_clk_stop_out_c3t ( stg4_mcu1_io_clk_stop_c3t  ),
	.stg4_mio_clk_stop_out_c3t ( stg4_mio_clk_stop_c3t  ),
	.stg4_mio_io2x_sync_en_out_c3t ( stg4_mio_io2x_sync_en_c3t  ),
	.stg4_ncu_clk_stop_out_c3b ( stg4_ncu_clk_stop_c3b  ),
	.stg4_ncu_io_clk_stop_out_c3b ( stg4_ncu_io_clk_stop_c3b  ),
	.stg4_peu_io_clk_stop_out_c3b ( stg4_peu_io_clk_stop_c3b  ),
	.stg4_sii_clk_stop_out_c3b ( stg4_sii_clk_stop_c3b  ),
	.stg4_sii_io_clk_stop_out_c3b ( stg4_sii_io_clk_stop_c3b  ),
	.stg4_spc0_clk_stop_out_c3t ( stg4_spc0_clk_stop_c3t  ),
//	.stg4_spc1_clk_stop_out_c2b ( stg4_spc1_clk_stop_c2b  ),
	.stg4_spc2_clk_stop_out_c3b ( stg4_spc2_clk_stop_c3b  ),
//	.stg4_spc5_clk_stop_out_c2b ( stg4_spc5_clk_stop_c2b  ),
	.stg2_mcu0_clk_stop_in_c2t ( stg2_mcu0_clk_stop_c1t ),// UNDRIVEN stg2_mcu0_clk_stop_in_c2t 
	.stg2_mcu1_clk_stop_in_c2t ( stg2_mcu1_clk_stop_c1t ),// UNDRIVEN stg2_mcu1_clk_stop_in_c2t 
	.stg3_mcu0_clk_stop_out_c2t ( stg3_mcu0_clk_stop_c2t ),
	.stg3_mcu1_clk_stop_out_c2t ( stg3_mcu1_clk_stop_c2t ),
  .cmp_gclk_c1_ccu(cmp_gclk_c1_ccu),
  .cmp_gclk_c2_ccx_left(cmp_gclk_c2_ccx_left),
  .cmp_gclk_c2_ccx_right(cmp_gclk_c2_ccx_right),
  .cmp_gclk_c3_db0(cmp_gclk_c3_db0),
  .cmp_gclk_c1_db1(cmp_gclk_c1_db1),
  .cmp_gclk_c3_dmu(cmp_gclk_c3_dmu),
  .cmp_gclk_c1_efu(cmp_gclk_c1_efu),
  .cmp_gclk_c3_l2b0(cmp_gclk_c3_l2b0),
  .cmp_gclk_c3_l2b1(cmp_gclk_c3_l2b1),
  .cmp_gclk_c3_l2b2(cmp_gclk_c3_l2b2),
  .cmp_gclk_c3_l2b3(cmp_gclk_c3_l2b3),
  .cmp_gclk_c1_l2b4(cmp_gclk_c1_l2b4),
  .cmp_gclk_c1_l2b5(cmp_gclk_c1_l2b5),
  .cmp_gclk_c1_l2b6(cmp_gclk_c1_l2b6),
  .cmp_gclk_c1_l2b7(cmp_gclk_c1_l2b7),
  .cmp_gclk_c3_l2d0(cmp_gclk_c3_l2d0),
  .cmp_gclk_c3_l2d1(cmp_gclk_c3_l2d1),
  .cmp_gclk_c3_l2d2(cmp_gclk_c3_l2d2),
  .cmp_gclk_c3_l2d3(cmp_gclk_c3_l2d3),
  .cmp_gclk_c1_l2d4(cmp_gclk_c1_l2d4),
  .cmp_gclk_c1_l2d5(cmp_gclk_c1_l2d5),
  .cmp_gclk_c1_l2d6(cmp_gclk_c1_l2d6),
  .cmp_gclk_c1_l2d7(cmp_gclk_c1_l2d7),
  .cmp_gclk_c3_l2t0(cmp_gclk_c3_l2t0),
  .cmp_gclk_c3_l2t2(cmp_gclk_c3_l2t2),
  .cmp_gclk_c1_l2t4(cmp_gclk_c1_l2t4),
  .cmp_gclk_c1_l2t6(cmp_gclk_c1_l2t6),
  .cmp_gclk_c2_l2t1(cmp_gclk_c2_l2t1),
  .cmp_gclk_c2_l2t3(cmp_gclk_c2_l2t3),
  .cmp_gclk_c2_l2t5(cmp_gclk_c2_l2t5),
  .cmp_gclk_c2_l2t7(cmp_gclk_c2_l2t7),
  .cmp_gclk_c4_mcu0(cmp_gclk_c4_mcu0),
  .cmp_gclk_c4_mcu1(cmp_gclk_c4_mcu1),
  .cmp_gclk_c0_mcu2(cmp_gclk_c0_mcu2),
  .cmp_gclk_c0_mcu3(cmp_gclk_c0_mcu3),
  .dr_gclk_c4_mcu0(dr_gclk_c4_mcu0),
  .dr_gclk_c4_mcu1(dr_gclk_c4_mcu1),
  .dr_gclk_c0_mcu2(dr_gclk_c0_mcu2),
  .dr_gclk_c0_mcu3(dr_gclk_c0_mcu3),
  .cmp_gclk_c1_mio(cmp_gclk_c1_mio),
  .cmp_gclk_c3_mio(cmp_gclk_c3_mio),
  .cmp_gclk_c2_mio_left(cmp_gclk_c2_mio_left),
  .cmp_gclk_c2_mio_right(cmp_gclk_c2_mio_right),
  .cmp_gclk_c3_ncu(cmp_gclk_c3_ncu),
  .cmp_gclk_c3_peu(cmp_gclk_c3_peu),
  .cmp_gclk_c3_sii(cmp_gclk_c3_sii),
  .cmp_gclk_c1_sio(cmp_gclk_c1_sio),
  .cmp_gclk_c3_spc0(cmp_gclk_c3_spc0),
  .cmp_gclk_c3_spc2(cmp_gclk_c3_spc2),
  .cmp_gclk_c1_spc4(cmp_gclk_c1_spc4),
  .cmp_gclk_c1_spc6(cmp_gclk_c1_spc6),
  .cmp_gclk_c2_spc1(cmp_gclk_c2_spc1),
  .cmp_gclk_c2_spc3(cmp_gclk_c2_spc3),
  .cmp_gclk_c2_spc5(cmp_gclk_c2_spc5),
  .cmp_gclk_c2_spc7(cmp_gclk_c2_spc7),
  .cmp_gclk_c1_tcu(cmp_gclk_c1_tcu),
  .cmp_gclk_c1_mac(cmp_gclk_c1_mac),
  .cmp_gclk_c0_rdp(cmp_gclk_c0_rdp),
  .cmp_gclk_c0_rtx(cmp_gclk_c0_rtx),
  .cmp_gclk_c0_tds(cmp_gclk_c0_tds),
  .cmp_gclk_c3_rng(cmp_gclk_c3_rng),
  .dr_gclk_c4_fsr0_0(dr_gclk_c4_fsr0_0),
  .dr_gclk_c4_fsr0_1(dr_gclk_c4_fsr0_1),
  .dr_gclk_c4_fsr0_2(dr_gclk_c4_fsr0_2),
  .dr_gclk_c4_fsr1_0(dr_gclk_c4_fsr1_0),
  .dr_gclk_c4_fsr1_1(dr_gclk_c4_fsr1_1),
  .dr_gclk_c4_fsr1_2(dr_gclk_c4_fsr1_2),
  .dr_gclk_c4_fsr2_0(dr_gclk_c4_fsr2_0),
  .dr_gclk_c4_fsr2_1(dr_gclk_c4_fsr2_1),
  .dr_gclk_c4_fsr2_2(dr_gclk_c4_fsr2_2),
  .dr_gclk_c4_fsr3_0(dr_gclk_c4_fsr3_0),
  .dr_gclk_c4_fsr3_1(dr_gclk_c4_fsr3_1),
  .dr_gclk_c4_fsr3_2(dr_gclk_c4_fsr3_2),
  .dr_gclk_c0_fsr4_0(dr_gclk_c0_fsr4_0),
  .dr_gclk_c0_fsr4_1(dr_gclk_c0_fsr4_1),
  .dr_gclk_c0_fsr4_2(dr_gclk_c0_fsr4_2),
  .dr_gclk_c0_fsr5_0(dr_gclk_c0_fsr5_0),
  .dr_gclk_c0_fsr5_1(dr_gclk_c0_fsr5_1),
  .dr_gclk_c0_fsr5_2(dr_gclk_c0_fsr5_2),
  .dr_gclk_c0_fsr6_0(dr_gclk_c0_fsr6_0),
  .dr_gclk_c0_fsr6_1(dr_gclk_c0_fsr6_1),
  .dr_gclk_c0_fsr6_2(dr_gclk_c0_fsr6_2),
  .dr_gclk_c2_fsr7_0(dr_gclk_c2_fsr7_0),
  .dr_gclk_c2_fsr7_1(dr_gclk_c2_fsr7_1),
  .dr_gclk_c2_fsr7_2(dr_gclk_c2_fsr7_2),
  .ccu_cmp_io_sync_en(ccu_cmp_io_sync_en),
  .ccu_dr_sync_en(ccu_dr_sync_en),
  .ccu_io2x_out(ccu_io2x_out),
  .ccu_io2x_sync_en(ccu_io2x_sync_en),
  .ccu_io_cmp_sync_en(ccu_io_cmp_sync_en),
  .ccu_io_out(ccu_io_out),
  .ccu_vco_aligned(ccu_vco_aligned),
  .gclk_aligned(gclk_aligned),
  .gl_ccu_clk_stop(gl_ccu_clk_stop),
  .gl_ccu_io_clk_stop(gl_ccu_io_clk_stop),
  .gl_ccx_clk_stop(gl_ccx_clk_stop),
  .gl_cmp_io_sync_en_c1b(gl_cmp_io_sync_en_c1b),
  .gl_cmp_io_sync_en_c1m(gl_cmp_io_sync_en_c1m),
  .gl_cmp_io_sync_en_c1t(gl_cmp_io_sync_en_c1t),
  .gl_cmp_io_sync_en_c2b(gl_cmp_io_sync_en_c2b),
  .gl_cmp_io_sync_en_c2t(gl_cmp_io_sync_en_c2t),
  .gl_cmp_io_sync_en_c3b(gl_cmp_io_sync_en_c3b),
  .gl_cmp_io_sync_en_c3t(gl_cmp_io_sync_en_c3t),
  .gl_cmp_io_sync_en_c3t0(gl_cmp_io_sync_en_c3t0),
  .gl_db0_clk_stop(gl_db0_clk_stop),
  .gl_db1_clk_stop(gl_db1_clk_stop),
  .gl_dmu_io_clk_stop(gl_dmu_io_clk_stop),
  .gl_dmu_peu_por_c3b(gl_dmu_peu_por_c3b),
  .gl_dmu_peu_wmr_c3b(gl_dmu_peu_wmr_c3b),
  .gl_dr_sync_en_c1m(gl_dr_sync_en_c1m),
  .gl_dr_sync_en_c3t(gl_dr_sync_en_c3t),
  .gl_efu_clk_stop(gl_efu_clk_stop),
  .gl_efu_io_clk_stop(gl_efu_io_clk_stop),
  .gl_io2x_out_c1b(gl_io2x_out_c1b),
  .gl_io2x_sync_en_c1m(gl_io2x_sync_en_c1m),
  .gl_io2x_sync_en_c3t(gl_io2x_sync_en_c3t),
  .gl_io2x_sync_en_c3t0(gl_io2x_sync_en_c3t0),
  .gl_io2x_sync_en_c2t(gl_io2x_sync_en_c2t),
  .gl_io_cmp_sync_en_c1b(gl_io_cmp_sync_en_c1b),
  .gl_io_cmp_sync_en_c1m(gl_io_cmp_sync_en_c1m),
  .gl_io_cmp_sync_en_c1t(gl_io_cmp_sync_en_c1t),
  .gl_io_cmp_sync_en_c2b(gl_io_cmp_sync_en_c2b),
  .gl_io_cmp_sync_en_c2t(gl_io_cmp_sync_en_c2t),
  .gl_io_cmp_sync_en_c3b(gl_io_cmp_sync_en_c3b),
  .gl_io_cmp_sync_en_c3t(gl_io_cmp_sync_en_c3t),
  .gl_io_cmp_sync_en_c3t0(gl_io_cmp_sync_en_c3t0),
  .gl_io_out_c1b(gl_io_out_c1b),
  .gl_io_out_c1m(gl_io_out_c1m),
  .gl_io_out_c3b(gl_io_out_c3b),
  .gl_io_out_c3b0(gl_io_out_c3b0),
  .gl_io_out_c3t(gl_io_out_c3t),
  .gl_l2_por_c1t(gl_l2_por_c1t),
  .gl_l2_por_c2b(gl_l2_por_c2b),
  .gl_l2_por_c2t(gl_l2_por_c2t),
  .gl_l2_por_c3b0(gl_l2_por_c3b0),
  .gl_l2_por_c3t(gl_l2_por_c3t),
  .gl_l2_por_c3t0(gl_l2_por_c3t0),
  .gl_l2_wmr_c1b(gl_l2_wmr_c1b),
  .gl_l2_wmr_c1t(gl_l2_wmr_c1t),
  .gl_l2_wmr_c2b(gl_l2_wmr_c2b),
  .gl_l2_wmr_c2t(gl_l2_wmr_c2t),
  .gl_l2_wmr_c3b(gl_l2_wmr_c3b),
  .gl_l2_wmr_c3t(gl_l2_wmr_c3t),
  .gl_l2_wmr_c3t0(gl_l2_wmr_c3t0),
  .gl_l2b0_clk_stop(gl_l2b0_clk_stop),
  .gl_l2b1_clk_stop(gl_l2b1_clk_stop),
  .gl_l2b2_clk_stop(gl_l2b2_clk_stop),
  .gl_l2b3_clk_stop(gl_l2b3_clk_stop),
  .gl_l2b4_clk_stop(gl_l2b4_clk_stop),
  .gl_l2b5_clk_stop(gl_l2b5_clk_stop),
  .gl_l2b6_clk_stop(gl_l2b6_clk_stop),
  .gl_l2b7_clk_stop(gl_l2b7_clk_stop),
  .gl_l2d0_clk_stop(gl_l2d0_clk_stop),
  .gl_l2d1_clk_stop(gl_l2d1_clk_stop),
  .gl_l2d2_clk_stop(gl_l2d2_clk_stop),
  .gl_l2d3_clk_stop(gl_l2d3_clk_stop),
  .gl_l2d4_clk_stop(gl_l2d4_clk_stop),
  .gl_l2d5_clk_stop(gl_l2d5_clk_stop),
  .gl_l2d6_clk_stop(gl_l2d6_clk_stop),
  .gl_l2d7_clk_stop(gl_l2d7_clk_stop),
  .gl_l2t0_clk_stop(gl_l2t0_clk_stop),
  .gl_l2t1_clk_stop(gl_l2t1_clk_stop),
  .gl_l2t2_clk_stop(gl_l2t2_clk_stop),
  .gl_l2t3_clk_stop(gl_l2t3_clk_stop),
  .gl_l2t4_clk_stop(gl_l2t4_clk_stop),
  .gl_l2t5_clk_stop(gl_l2t5_clk_stop),
  .gl_l2t6_clk_stop(gl_l2t6_clk_stop),
  .gl_l2t7_clk_stop(gl_l2t7_clk_stop),
  .gl_mac_io_clk_stop(gl_mac_io_clk_stop),
  .gl_mcu0_clk_stop(gl_mcu0_clk_stop),
  .gl_mcu0_dr_clk_stop(gl_mcu0_dr_clk_stop),
  .gl_mcu0_io_clk_stop(gl_mcu0_io_clk_stop),
  .gl_mcu1_clk_stop(gl_mcu1_clk_stop),
  .gl_mcu1_dr_clk_stop(gl_mcu1_dr_clk_stop),
  .gl_mcu1_io_clk_stop(gl_mcu1_io_clk_stop),
  .gl_mcu2_clk_stop(gl_mcu2_clk_stop),
  .gl_mcu2_dr_clk_stop(gl_mcu2_dr_clk_stop),
  .gl_mcu2_io_clk_stop(gl_mcu2_io_clk_stop),
  .gl_mcu3_clk_stop(gl_mcu3_clk_stop),
  .gl_mcu3_dr_clk_stop(gl_mcu3_dr_clk_stop),
  .gl_mcu3_io_clk_stop(gl_mcu3_io_clk_stop),
  .gl_mio_clk_stop_c1t(gl_mio_clk_stop_c1t),
  .gl_mio_clk_stop_c2t(gl_mio_clk_stop_c2t),
  .gl_mio_clk_stop_c3t(gl_mio_clk_stop_c3t),
  .gl_mio_io2x_sync_en_c1t(gl_mio_io2x_sync_en_c1t),
  .gl_ncu_clk_stop(gl_ncu_clk_stop),
  .gl_ncu_io_clk_stop(gl_ncu_io_clk_stop),
  .gl_peu_io_clk_stop(gl_peu_io_clk_stop),
  .gl_rdp_io_clk_stop(gl_rdp_io_clk_stop),
  .gl_rst_clk_stop(gl_rst_clk_stop),
  .gl_rst_io_clk_stop(gl_rst_io_clk_stop),
  .gl_rst_l2_por_c1m(gl_rst_l2_por_c1m),
  .gl_rst_l2_wmr_c1m(gl_rst_l2_wmr_c1m),
  .gl_rst_mac_c1b(gl_rst_mac_c1b),
  .gl_rst_niu_wmr_c1b(gl_rst_niu_wmr_c1b),
  .gl_rtx_io_clk_stop(gl_rtx_io_clk_stop),
  .gl_sii_clk_stop(gl_sii_clk_stop),
  .gl_sii_io_clk_stop(gl_sii_io_clk_stop),
  .gl_sio_clk_stop(gl_sio_clk_stop),
  .gl_sio_io_clk_stop(gl_sio_io_clk_stop),
  .gl_spc0_clk_stop(gl_spc0_clk_stop),
  .gl_spc1_clk_stop(gl_spc1_clk_stop),
  .gl_spc2_clk_stop(gl_spc2_clk_stop),
  .gl_spc3_clk_stop(gl_spc3_clk_stop),
  .gl_spc4_clk_stop(gl_spc4_clk_stop),
  .gl_spc5_clk_stop(gl_spc5_clk_stop),
  .gl_spc6_clk_stop(gl_spc6_clk_stop),
  .gl_spc7_clk_stop(gl_spc7_clk_stop),
  .gl_tds_io_clk_stop(gl_tds_io_clk_stop),
  .rst_dmu_peu_por_(rst_dmu_peu_por_),
  .rst_dmu_peu_wmr_(rst_dmu_peu_wmr_),
  .rst_l2_por_(rst_l2_por_),
  .rst_l2_wmr_(rst_l2_wmr_),
  .rst_niu_mac_(rst_niu_mac_),
  .gl_l2_por_c1b(gl_l2_por_c1b),
  .rst_niu_wmr_(rst_niu_wmr_),
  .tcu_ccu_clk_stop(tcu_ccu_clk_stop),
  .tcu_ccu_io_clk_stop(tcu_ccu_io_clk_stop),
  .tcu_ccx_clk_stop(tcu_ccx_clk_stop),
  .tcu_db0_clk_stop(tcu_db0_clk_stop),
  .tcu_db1_clk_stop(tcu_db1_clk_stop),
  .tcu_dmu_io_clk_stop(tcu_dmu_io_clk_stop),
  .tcu_efu_clk_stop(tcu_efu_clk_stop),
  .tcu_efu_io_clk_stop(tcu_efu_io_clk_stop),
  .tcu_l2b0_clk_stop(tcu_l2b0_clk_stop),
  .tcu_l2b1_clk_stop(tcu_l2b1_clk_stop),
  .tcu_l2b2_clk_stop(tcu_l2b2_clk_stop),
  .tcu_l2b3_clk_stop(tcu_l2b3_clk_stop),
  .tcu_l2b4_clk_stop(tcu_l2b4_clk_stop),
  .tcu_l2b5_clk_stop(tcu_l2b5_clk_stop),
  .tcu_l2b6_clk_stop(tcu_l2b6_clk_stop),
  .tcu_l2b7_clk_stop(tcu_l2b7_clk_stop),
  .tcu_l2d0_clk_stop(tcu_l2d0_clk_stop),
  .tcu_l2d1_clk_stop(tcu_l2d1_clk_stop),
  .tcu_l2d2_clk_stop(tcu_l2d2_clk_stop),
  .tcu_l2d3_clk_stop(tcu_l2d3_clk_stop),
  .tcu_l2d4_clk_stop(tcu_l2d4_clk_stop),
  .tcu_l2d5_clk_stop(tcu_l2d5_clk_stop),
  .tcu_l2d6_clk_stop(tcu_l2d6_clk_stop),
  .tcu_l2d7_clk_stop(tcu_l2d7_clk_stop),
  .tcu_l2t0_clk_stop(tcu_l2t0_clk_stop),
  .tcu_l2t1_clk_stop(tcu_l2t1_clk_stop),
  .tcu_l2t2_clk_stop(tcu_l2t2_clk_stop),
  .tcu_l2t3_clk_stop(tcu_l2t3_clk_stop),
  .tcu_l2t4_clk_stop(tcu_l2t4_clk_stop),
  .tcu_l2t5_clk_stop(tcu_l2t5_clk_stop),
  .tcu_l2t6_clk_stop(tcu_l2t6_clk_stop),
  .tcu_l2t7_clk_stop(tcu_l2t7_clk_stop),
  .tcu_mac_io_clk_stop(tcu_mac_io_clk_stop),
  .tcu_mcu0_clk_stop(tcu_mcu0_clk_stop),
  .tcu_mcu0_dr_clk_stop(tcu_mcu0_dr_clk_stop),
  .tcu_mcu0_io_clk_stop(tcu_mcu0_io_clk_stop),
  .tcu_mcu1_clk_stop(tcu_mcu1_clk_stop),
  .tcu_mcu1_dr_clk_stop(tcu_mcu1_dr_clk_stop),
  .tcu_mcu1_io_clk_stop(tcu_mcu1_io_clk_stop),
  .tcu_mcu2_clk_stop(tcu_mcu2_clk_stop),
  .tcu_mcu2_dr_clk_stop(tcu_mcu2_dr_clk_stop),
  .tcu_mcu2_io_clk_stop(tcu_mcu2_io_clk_stop),
  .tcu_mcu3_clk_stop(tcu_mcu3_clk_stop),
  .tcu_mcu3_dr_clk_stop(tcu_mcu3_dr_clk_stop),
  .tcu_mcu3_io_clk_stop(tcu_mcu3_io_clk_stop),
  .tcu_mio_clk_stop(tcu_mio_clk_stop),
  .tcu_ncu_clk_stop(tcu_ncu_clk_stop),
  .tcu_ncu_io_clk_stop(tcu_ncu_io_clk_stop),
  .tcu_peu_io_clk_stop(tcu_peu_io_clk_stop),
  .tcu_rdp_io_clk_stop(tcu_rdp_io_clk_stop),
  .tcu_rst_clk_stop(tcu_rst_clk_stop),
  .tcu_rst_io_clk_stop(tcu_rst_io_clk_stop),
  .tcu_rtx_io_clk_stop(tcu_rtx_io_clk_stop),
  .tcu_sii_clk_stop(tcu_sii_clk_stop),
  .tcu_sii_io_clk_stop(tcu_sii_io_clk_stop),
  .tcu_sio_clk_stop(tcu_sio_clk_stop),
  .tcu_sio_io_clk_stop(tcu_sio_io_clk_stop),
  .tcu_spc0_clk_stop(tcu_spc0_clk_stop),
  .tcu_spc1_clk_stop(tcu_spc1_clk_stop),
  .tcu_spc2_clk_stop(tcu_spc2_clk_stop),
  .tcu_spc3_clk_stop(tcu_spc3_clk_stop),
  .tcu_spc4_clk_stop(tcu_spc4_clk_stop),
  .tcu_spc5_clk_stop(tcu_spc5_clk_stop),
  .tcu_spc6_clk_stop(tcu_spc6_clk_stop),
  .tcu_spc7_clk_stop(tcu_spc7_clk_stop),
  .tcu_tds_io_clk_stop(tcu_tds_io_clk_stop)
    // PRIMARY OUTPUTS (CLKS) -- AUTOMATIC CONNECTIONS
	// PRIMARY OUTPUTS -- AUTOMATIC CONNECTIONS
);



endmodule // cpu


