// Small test module

module sub_and (
input wire d,
input wire b,
output wire out);

assign out = d & b;

endmodule
