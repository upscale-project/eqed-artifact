module xtest_checker_bind;

   bind xtest xtest_checker check1 (.a_ch(a),.clk(clk));

endmodule // xtest_checker_bind

   