module inst_constraint_bind;

   bind spc_wrapper.spc.dec inst_constraint inst_constraint_0 (.clk(l2clk),
                                                               .dec_valid_d(dec_valid0_d),
                                                               .instruction(ifu_buf0_inst0));

endmodule // inst_constraint_bind



   
