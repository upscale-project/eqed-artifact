`include "qed.vh"


module l2c_checker2 (/*AUTOARG*/
   // Inputs
   clk, rst, ena  
   );

   input        clk;
   input        rst;
   input        ena;
    
   genvar       j;




   
   // PROPERTIES
   

   // ASSUMPTIONS
   



   // ASSERTIONS



endmodule // l2c_checker2
