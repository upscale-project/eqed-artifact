
module dff3 (
input [2:0] d,
output wire [2:0] q);

assign q = d*2;

endmodule
