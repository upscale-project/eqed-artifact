// test dff module - just for parsing (nto the real dff module)
// functionality does not work

module dff (input d,
            input clk,
	    output q);

assign q = d;

endmodule
