/* small test submodule */

module add
(
input wire d,
input wire b_add,
output wire out_add
);

assign out_add = d + b_add;

endmodule
